* SPICE3 file created from multiplier_test.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY=5
.option scale=0.09u
.global vdd gnd


Vdd vdd gnd 'SUPPLY'

* Inputs for testing the functionality
vinA0 inA0 gnd pulse 0 'SUPPLY' 0ns 0.1ns 0.1ns 10ns 20ns
vinA1 inA1 gnd pulse 0 'SUPPLY' 10ns 0.1ns 0.1ns 10ns 20ns
vinA2 inA2 gnd pulse 0 'SUPPLY' 10ns 0.1ns 0.1ns 10ns 20ns
vinA3 inA3 gnd pulse 0 'SUPPLY' 0ns 0.1ns 0.1ns 10ns 20ns

vinB0 inB0 gnd pulse 0 'SUPPLY' 0ns 0.1ns 0.1ns 20ns 40ns
vinB1 inB1 gnd pulse 0 'SUPPLY' 10ns 0.1ns 0.1ns 20ns 40ns
vinB2 inB2 gnd pulse 0 'SUPPLY' 0ns 0.1ns 0.1ns 20ns 40ns
vinB3 inB3 gnd pulse 0 'SUPPLY' 0ns 0.1ns 0.1ns 20ns 40ns
* vinC inC gnd pulse 0 'SUPPLY' 0ns 0.1ns 0.1ns 40ns 80ns

* Inputs for calculating Delays
* va inA0 gnd 'SUPPLY' DC
* vb inA1 gnd 0 DC
* vc inA2 gnd pulse 'SUPPLY' 0 0ns 10ps 10ps 10ns 20ns
* vd inA3 gnd 'SUPPLY' DC

* ve inB0 gnd pulse 0 'SUPPLY' 0ns 10ps 10ps 10ns 20ns
* vf inB1 gnd pulse 0 'SUPPLY' 0ns 10ps 10ps 10ns 20ns
* vg inB2 gnd pulse 'SUPPLY' 0 0ns 10ps 10ps 10ns 20ns
* vh inB3 gnd 'SUPPLY' DC

* vinA0 inA0 gnd 1 DC
* vinA1 inA1 gnd 1 DC
* vinA2 inA2 gnd 1 DC
* vinA3 inA3 gnd 1 DC

* vinB0 inB0 gnd 1 DC
* vinB1 inB1 gnd 1 DC
* vinB2 inB2 gnd 1 DC
* vinB3 inB3 gnd 1 DC



M1000 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n611_n78# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1001 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n2157_n115# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=13580 ps=6190
M1002 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n611_n78# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=15840 ps=6850
M1003 vdd multiplier_0/m1_n2157_n115# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1004 multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1005 multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1006 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1007 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n2157_n115# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1008 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1009 vdd multiplier_0/m1_n2157_n115# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1010 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n611_n78# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1011 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n2157_n115# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1012 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n611_n78# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1013 vdd multiplier_0/m1_n2157_n115# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1014 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n611_n78# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1015 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1016 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n611_n78# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1017 vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1018 multiplier_0/4bitadder_0/fulladder_0/m1_411_129# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1019 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1020 multiplier_0/4bitadder_0/fulladder_0/m1_411_129# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1021 vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1022 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/m1_n594_383# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1023 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1024 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/m1_n594_383# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1025 vdd multiplier_0/4bitadder_0/fulladder_0/m1_411_129# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1026 multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1027 multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1028 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1029 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1030 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1031 vdd multiplier_0/4bitadder_0/fulladder_0/m1_411_129# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1032 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/m1_n594_383# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1033 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1034 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/m1_n594_383# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1035 vdd multiplier_0/4bitadder_0/fulladder_0/m1_411_129# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1036 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/m1_n594_383# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1037 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1038 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/m1_n594_383# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1039 vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1040 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1041 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1042 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1043 vdd multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1044 multiplier_0/4bitadder_0/m1_n1726_385# multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1045 multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1046 multiplier_0/4bitadder_0/m1_n1726_385# multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# vdd multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1047 vdd multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_0/m1_n1726_385# multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1048 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1049 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# vdd multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1050 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1051 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# vdd multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_1/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1052 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n980_n67# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1053 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n2469_n98# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1054 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n980_n67# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1055 vdd multiplier_0/m1_n2469_n98# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1056 multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1057 multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1058 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1059 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n2469_n98# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1060 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1061 vdd multiplier_0/m1_n2469_n98# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1062 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n980_n67# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1063 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n2469_n98# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1064 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n980_n67# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1065 vdd multiplier_0/m1_n2469_n98# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1066 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n980_n67# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1067 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1068 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n980_n67# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1069 vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1070 multiplier_0/4bitadder_0/fulladder_1/m1_411_129# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1071 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1072 multiplier_0/4bitadder_0/fulladder_1/m1_411_129# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1073 vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_1/m1_411_129# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1074 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/m1_n1726_385# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1075 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/fulladder_1/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1076 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/m1_n1726_385# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1077 vdd multiplier_0/4bitadder_0/fulladder_1/m1_411_129# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1078 multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1079 multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1080 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1081 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# multiplier_0/4bitadder_0/fulladder_1/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1082 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1083 vdd multiplier_0/4bitadder_0/fulladder_1/m1_411_129# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1084 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/m1_n1726_385# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1085 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/fulladder_1/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1086 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/m1_n1726_385# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1087 vdd multiplier_0/4bitadder_0/fulladder_1/m1_411_129# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1088 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/m1_n1726_385# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1089 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1090 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/m1_n1726_385# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1091 vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1092 multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1093 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1094 multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1095 vdd multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1096 multiplier_0/4bitadder_0/m1_n2858_385# multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1097 multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1098 multiplier_0/4bitadder_0/m1_n2858_385# multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# vdd multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1099 vdd multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_0/m1_n2858_385# multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1100 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1101 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# vdd multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1102 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1103 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# vdd multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_1/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1104 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# gnd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1105 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n2782_n115# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1106 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# gnd vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1107 vdd multiplier_0/m1_n2782_n115# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1108 multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1109 multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1110 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1111 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n2782_n115# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1112 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1113 vdd multiplier_0/m1_n2782_n115# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1114 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# gnd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1115 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n2782_n115# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1116 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# gnd vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1117 vdd multiplier_0/m1_n2782_n115# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1118 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# gnd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1119 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1120 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# gnd vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1121 vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1122 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1123 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1124 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1125 vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1126 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/m1_n2858_385# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1127 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/fulladder_2/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1128 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/m1_n2858_385# vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1129 vdd multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1130 multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1131 multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1132 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1133 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# multiplier_0/4bitadder_0/fulladder_2/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1134 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1135 vdd multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1136 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/m1_n2858_385# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1137 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/fulladder_2/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1138 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/m1_n2858_385# vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1139 vdd multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1140 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/m1_n2858_385# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1141 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1142 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/m1_n2858_385# vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1143 vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1144 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1145 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1146 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1147 vdd multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1148 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1149 multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1150 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# vdd multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1151 vdd multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1152 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1153 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# vdd multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1154 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1155 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# vdd multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_1/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1156 multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n294_n107# multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1157 multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n1820_n104# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1158 multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n294_n107# vdd multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1159 vdd multiplier_0/m1_n1820_n104# multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1160 multiplier_0/4bitadder_0/m1_n594_383# multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1161 multiplier_0/4bitadder_0/m1_n594_383# multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_0/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1162 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1163 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n1820_n104# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1164 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1165 vdd multiplier_0/m1_n1820_n104# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1166 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n294_n107# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1167 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n1820_n104# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1168 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n294_n107# vdd multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1169 vdd multiplier_0/m1_n1820_n104# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1170 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n294_n107# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1171 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1172 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n294_n107# vdd multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1173 vdd multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1174 P1 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1175 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1176 P1 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1177 vdd multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# P1 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1178 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1179 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n2968_n1347# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1180 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n1473_n1361# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1181 vdd multiplier_0/m1_n2968_n1347# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1182 multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1183 multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1184 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1185 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n2968_n1347# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1186 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1187 vdd multiplier_0/m1_n2968_n1347# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1188 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1189 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n2968_n1347# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1190 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n1473_n1361# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1191 vdd multiplier_0/m1_n2968_n1347# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1192 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1193 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1194 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n1473_n1361# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1195 vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1196 multiplier_0/4bitadder_1/fulladder_0/m1_411_129# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1197 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1198 multiplier_0/4bitadder_1/fulladder_0/m1_411_129# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1199 vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1200 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/m1_n594_383# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1201 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1202 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/m1_n594_383# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1203 vdd multiplier_0/4bitadder_1/fulladder_0/m1_411_129# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1204 multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1205 multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1206 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1207 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1208 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1209 vdd multiplier_0/4bitadder_1/fulladder_0/m1_411_129# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1210 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/m1_n594_383# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1211 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1212 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/m1_n594_383# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1213 vdd multiplier_0/4bitadder_1/fulladder_0/m1_411_129# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1214 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/m1_n594_383# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1215 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1216 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/m1_n594_383# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1217 vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1218 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1219 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1220 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1221 vdd multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1222 multiplier_0/4bitadder_1/m1_n1726_385# multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1223 multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1224 multiplier_0/4bitadder_1/m1_n1726_385# multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# vdd multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1225 vdd multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_1/m1_n1726_385# multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1226 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1227 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# vdd multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1228 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1229 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# vdd multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_1/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1230 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1231 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n3306_n1348# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1232 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2288_n756# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1233 vdd multiplier_0/m1_n3306_n1348# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1234 multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1235 multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1236 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1237 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n3306_n1348# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1238 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1239 vdd multiplier_0/m1_n3306_n1348# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1240 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1241 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n3306_n1348# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1242 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2288_n756# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1243 vdd multiplier_0/m1_n3306_n1348# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1244 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1245 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1246 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n2288_n756# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1247 vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1248 multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1249 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1250 multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1251 vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1252 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/m1_n1726_385# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1253 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/fulladder_1/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1254 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/m1_n1726_385# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1255 vdd multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1256 multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1257 multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1258 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1259 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# multiplier_0/4bitadder_1/fulladder_1/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1260 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1261 vdd multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1262 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/m1_n1726_385# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1263 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/fulladder_1/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1264 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/m1_n1726_385# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1265 vdd multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1266 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/m1_n1726_385# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1267 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1268 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/m1_n1726_385# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1269 vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1270 multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1271 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1272 multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1273 vdd multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1274 multiplier_0/4bitadder_1/m1_n2858_385# multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1275 multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1276 multiplier_0/4bitadder_1/m1_n2858_385# multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# vdd multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1277 vdd multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_1/m1_n2858_385# multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1278 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1279 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# vdd multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1280 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1281 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# vdd multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_1/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1282 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1283 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n3602_n1349# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1284 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n3416_n801# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1285 vdd multiplier_0/m1_n3602_n1349# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1286 multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1287 multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1288 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1289 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n3602_n1349# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1290 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1291 vdd multiplier_0/m1_n3602_n1349# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1292 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1293 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n3602_n1349# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1294 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n3416_n801# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1295 vdd multiplier_0/m1_n3602_n1349# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1296 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1297 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1298 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n3416_n801# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1299 vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1300 multiplier_0/4bitadder_1/fulladder_2/m1_411_129# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1301 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1302 multiplier_0/4bitadder_1/fulladder_2/m1_411_129# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1303 vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_2/m1_411_129# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1304 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/m1_n2858_385# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1305 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/fulladder_2/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1306 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/m1_n2858_385# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1307 vdd multiplier_0/4bitadder_1/fulladder_2/m1_411_129# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1308 multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1309 multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1310 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1311 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# multiplier_0/4bitadder_1/fulladder_2/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1312 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1313 vdd multiplier_0/4bitadder_1/fulladder_2/m1_411_129# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1314 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/m1_n2858_385# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1315 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/fulladder_2/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1316 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/m1_n2858_385# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1317 vdd multiplier_0/4bitadder_1/fulladder_2/m1_411_129# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1318 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/m1_n2858_385# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1319 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1320 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/m1_n2858_385# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1321 vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1322 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1323 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1324 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1325 vdd multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1326 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1327 multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1328 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# vdd multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1329 vdd multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1330 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1331 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# vdd multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1332 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1333 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# vdd multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_1/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1334 multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1335 multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n2617_n1342# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1336 multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n1128_n767# vdd multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1337 vdd multiplier_0/m1_n2617_n1342# multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1338 multiplier_0/4bitadder_1/m1_n594_383# multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1339 multiplier_0/4bitadder_1/m1_n594_383# multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_1/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1340 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1341 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n2617_n1342# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1342 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1343 vdd multiplier_0/m1_n2617_n1342# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1344 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1345 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n2617_n1342# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1346 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n1128_n767# vdd multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1347 vdd multiplier_0/m1_n2617_n1342# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1348 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1349 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1350 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n1128_n767# vdd multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1351 vdd multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1352 P2 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1353 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1354 P2 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1355 vdd multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# P2 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1356 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1357 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n4201_n2800# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1358 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2688_n2050# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1359 vdd multiplier_0/m1_n4201_n2800# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1360 multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1361 multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1362 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1363 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n4201_n2800# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1364 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1365 vdd multiplier_0/m1_n4201_n2800# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1366 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1367 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n4201_n2800# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1368 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2688_n2050# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1369 vdd multiplier_0/m1_n4201_n2800# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1370 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1371 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1372 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n2688_n2050# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1373 vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1374 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1375 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1376 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1377 vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1378 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/m1_n594_383# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1379 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/fulladder_0/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1380 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/m1_n594_383# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1381 vdd multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1382 multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1383 multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1384 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1385 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# multiplier_0/4bitadder_2/fulladder_0/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1386 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1387 vdd multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1388 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/m1_n594_383# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1389 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/fulladder_0/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1390 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/m1_n594_383# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1391 vdd multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1392 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/m1_n594_383# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1393 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1394 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/m1_n594_383# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1395 vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1396 P4 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1397 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1398 P4 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1399 vdd multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# P4 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1400 multiplier_0/4bitadder_2/m1_n1726_385# multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1401 multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1402 multiplier_0/4bitadder_2/m1_n1726_385# multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# vdd multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1403 vdd multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_2/m1_n1726_385# multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1404 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1405 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# vdd multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1406 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1407 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# vdd multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_1/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1408 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1409 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n4533_n2563# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1410 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n3123_n2056# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1411 vdd multiplier_0/m1_n4533_n2563# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1412 multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1413 multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1414 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1415 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n4533_n2563# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1416 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1417 vdd multiplier_0/m1_n4533_n2563# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1418 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1419 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n4533_n2563# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1420 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n3123_n2056# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1421 vdd multiplier_0/m1_n4533_n2563# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1422 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1423 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1424 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n3123_n2056# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1425 vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1426 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1427 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1428 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1429 vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1430 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/m1_n1726_385# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1431 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/fulladder_1/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1432 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/m1_n1726_385# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1433 vdd multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1434 multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1435 multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1436 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1437 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# multiplier_0/4bitadder_2/fulladder_1/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1438 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1439 vdd multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1440 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/m1_n1726_385# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1441 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/fulladder_1/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1442 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/m1_n1726_385# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1443 vdd multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1444 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/m1_n1726_385# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1445 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1446 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/m1_n1726_385# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1447 vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1448 P5 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1449 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1450 P5 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1451 vdd multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# P5 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1452 multiplier_0/4bitadder_2/m1_n2858_385# multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1453 multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1454 multiplier_0/4bitadder_2/m1_n2858_385# multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# vdd multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1455 vdd multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_2/m1_n2858_385# multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1456 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1457 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# vdd multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1458 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1459 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# vdd multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_1/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1460 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1461 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n4992_n2575# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1462 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n4235_n2059# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1463 vdd multiplier_0/m1_n4992_n2575# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1464 multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1465 multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1466 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1467 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n4992_n2575# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1468 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1469 vdd multiplier_0/m1_n4992_n2575# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1470 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1471 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n4992_n2575# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1472 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n4235_n2059# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1473 vdd multiplier_0/m1_n4992_n2575# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1474 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1475 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1476 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n4235_n2059# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1477 vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1478 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1479 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1480 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1481 vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1482 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/m1_n2858_385# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1483 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/fulladder_2/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1484 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/m1_n2858_385# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1485 vdd multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1486 multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1487 multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1488 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1489 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# multiplier_0/4bitadder_2/fulladder_2/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1490 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1491 vdd multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1492 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/m1_n2858_385# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1493 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/fulladder_2/m1_411_129# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1494 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/m1_n2858_385# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1495 vdd multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1496 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/m1_n2858_385# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1497 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1498 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/m1_n2858_385# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1499 vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1500 P6 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1501 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1502 P6 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1503 vdd multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# P6 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1504 P7 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1505 multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1506 P7 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# vdd multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1507 vdd multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# P7 multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1508 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1509 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# vdd multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1510 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1511 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# vdd multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_1/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1512 multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1513 multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n3849_n2792# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1514 multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2369_n2126# vdd multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1515 vdd multiplier_0/m1_n3849_n2792# multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1516 multiplier_0/4bitadder_2/m1_n594_383# multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1517 multiplier_0/4bitadder_2/m1_n594_383# multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# vdd multiplier_0/4bitadder_2/halfadder_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1518 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1519 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/m1_n3849_n2792# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1520 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# vdd multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1521 vdd multiplier_0/m1_n3849_n2792# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1522 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1523 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n3849_n2792# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1524 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2369_n2126# vdd multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1525 vdd multiplier_0/m1_n3849_n2792# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1526 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1527 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1528 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n2369_n2126# vdd multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1529 vdd multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1530 P3 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1531 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/a_n5_n50# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1532 P3 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# vdd multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1533 vdd multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# P3 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1534 multiplier_0/and_0/m1_59_58# inA0 multiplier_0/and_0/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1535 multiplier_0/and_0/nand_0/a_n5_n50# inB0 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1536 multiplier_0/and_0/m1_59_58# inA0 vdd multiplier_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1537 vdd inB0 multiplier_0/and_0/m1_59_58# multiplier_0/and_0/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1538 P0 multiplier_0/and_0/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1539 P0 multiplier_0/and_0/m1_59_58# vdd multiplier_0/and_0/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1540 multiplier_0/and_1/m1_59_58# inA1 multiplier_0/and_1/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1541 multiplier_0/and_1/nand_0/a_n5_n50# inB0 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1542 multiplier_0/and_1/m1_59_58# inA1 vdd multiplier_0/and_1/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1543 vdd inB0 multiplier_0/and_1/m1_59_58# multiplier_0/and_1/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1544 multiplier_0/m1_n294_n107# multiplier_0/and_1/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1545 multiplier_0/m1_n294_n107# multiplier_0/and_1/m1_59_58# vdd multiplier_0/and_1/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1546 multiplier_0/and_2/m1_59_58# inA2 multiplier_0/and_2/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1547 multiplier_0/and_2/nand_0/a_n5_n50# inB0 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1548 multiplier_0/and_2/m1_59_58# inA2 vdd multiplier_0/and_2/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1549 vdd inB0 multiplier_0/and_2/m1_59_58# multiplier_0/and_2/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1550 multiplier_0/m1_n611_n78# multiplier_0/and_2/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1551 multiplier_0/m1_n611_n78# multiplier_0/and_2/m1_59_58# vdd multiplier_0/and_2/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1552 multiplier_0/and_3/m1_59_58# inA3 multiplier_0/and_3/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1553 multiplier_0/and_3/nand_0/a_n5_n50# inB0 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1554 multiplier_0/and_3/m1_59_58# inA3 vdd multiplier_0/and_3/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1555 vdd inB0 multiplier_0/and_3/m1_59_58# multiplier_0/and_3/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1556 multiplier_0/m1_n980_n67# multiplier_0/and_3/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1557 multiplier_0/m1_n980_n67# multiplier_0/and_3/m1_59_58# vdd multiplier_0/and_3/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1558 multiplier_0/and_4/m1_59_58# inA0 multiplier_0/and_4/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1559 multiplier_0/and_4/nand_0/a_n5_n50# inB1 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1560 multiplier_0/and_4/m1_59_58# inA0 vdd multiplier_0/and_4/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1561 vdd inB1 multiplier_0/and_4/m1_59_58# multiplier_0/and_4/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1562 multiplier_0/m1_n1820_n104# multiplier_0/and_4/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1563 multiplier_0/m1_n1820_n104# multiplier_0/and_4/m1_59_58# vdd multiplier_0/and_4/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1564 multiplier_0/and_5/m1_59_58# inA1 multiplier_0/and_5/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1565 multiplier_0/and_5/nand_0/a_n5_n50# inB1 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1566 multiplier_0/and_5/m1_59_58# inA1 vdd multiplier_0/and_5/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1567 vdd inB1 multiplier_0/and_5/m1_59_58# multiplier_0/and_5/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1568 multiplier_0/m1_n2157_n115# multiplier_0/and_5/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1569 multiplier_0/m1_n2157_n115# multiplier_0/and_5/m1_59_58# vdd multiplier_0/and_5/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1570 multiplier_0/and_6/m1_59_58# inA2 multiplier_0/and_6/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1571 multiplier_0/and_6/nand_0/a_n5_n50# inB1 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1572 multiplier_0/and_6/m1_59_58# inA2 vdd multiplier_0/and_6/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1573 vdd inB1 multiplier_0/and_6/m1_59_58# multiplier_0/and_6/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1574 multiplier_0/m1_n2469_n98# multiplier_0/and_6/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1575 multiplier_0/m1_n2469_n98# multiplier_0/and_6/m1_59_58# vdd multiplier_0/and_6/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1576 multiplier_0/and_7/m1_59_58# inA3 multiplier_0/and_7/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1577 multiplier_0/and_7/nand_0/a_n5_n50# inB1 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1578 multiplier_0/and_7/m1_59_58# inA3 vdd multiplier_0/and_7/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1579 vdd inB1 multiplier_0/and_7/m1_59_58# multiplier_0/and_7/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1580 multiplier_0/m1_n2782_n115# multiplier_0/and_7/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1581 multiplier_0/m1_n2782_n115# multiplier_0/and_7/m1_59_58# vdd multiplier_0/and_7/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1582 multiplier_0/and_8/m1_59_58# inA0 multiplier_0/and_8/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1583 multiplier_0/and_8/nand_0/a_n5_n50# inB2 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1584 multiplier_0/and_8/m1_59_58# inA0 vdd multiplier_0/and_8/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1585 vdd inB2 multiplier_0/and_8/m1_59_58# multiplier_0/and_8/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1586 multiplier_0/m1_n2617_n1342# multiplier_0/and_8/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1587 multiplier_0/m1_n2617_n1342# multiplier_0/and_8/m1_59_58# vdd multiplier_0/and_8/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1588 multiplier_0/and_9/m1_59_58# inA1 multiplier_0/and_9/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1589 multiplier_0/and_9/nand_0/a_n5_n50# inB2 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1590 multiplier_0/and_9/m1_59_58# inA1 vdd multiplier_0/and_9/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1591 vdd inB2 multiplier_0/and_9/m1_59_58# multiplier_0/and_9/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1592 multiplier_0/m1_n2968_n1347# multiplier_0/and_9/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1593 multiplier_0/m1_n2968_n1347# multiplier_0/and_9/m1_59_58# vdd multiplier_0/and_9/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1594 multiplier_0/and_10/m1_59_58# inA2 multiplier_0/and_10/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1595 multiplier_0/and_10/nand_0/a_n5_n50# inB2 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1596 multiplier_0/and_10/m1_59_58# inA2 vdd multiplier_0/and_10/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1597 vdd inB2 multiplier_0/and_10/m1_59_58# multiplier_0/and_10/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1598 multiplier_0/m1_n3306_n1348# multiplier_0/and_10/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1599 multiplier_0/m1_n3306_n1348# multiplier_0/and_10/m1_59_58# vdd multiplier_0/and_10/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1600 multiplier_0/and_11/m1_59_58# inA3 multiplier_0/and_11/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1601 multiplier_0/and_11/nand_0/a_n5_n50# inB2 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1602 multiplier_0/and_11/m1_59_58# inA3 vdd multiplier_0/and_11/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1603 vdd inB2 multiplier_0/and_11/m1_59_58# multiplier_0/and_11/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1604 multiplier_0/m1_n3602_n1349# multiplier_0/and_11/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1605 multiplier_0/m1_n3602_n1349# multiplier_0/and_11/m1_59_58# vdd multiplier_0/and_11/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1606 multiplier_0/and_12/m1_59_58# inA3 multiplier_0/and_12/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1607 multiplier_0/and_12/nand_0/a_n5_n50# inB3 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1608 multiplier_0/and_12/m1_59_58# inA3 vdd multiplier_0/and_12/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1609 vdd inB3 multiplier_0/and_12/m1_59_58# multiplier_0/and_12/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1610 multiplier_0/m1_n4992_n2575# multiplier_0/and_12/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1611 multiplier_0/m1_n4992_n2575# multiplier_0/and_12/m1_59_58# vdd multiplier_0/and_12/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1612 multiplier_0/and_13/m1_59_58# inA2 multiplier_0/and_13/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1613 multiplier_0/and_13/nand_0/a_n5_n50# inB3 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1614 multiplier_0/and_13/m1_59_58# inA2 vdd multiplier_0/and_13/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1615 vdd inB3 multiplier_0/and_13/m1_59_58# multiplier_0/and_13/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1616 multiplier_0/m1_n4533_n2563# multiplier_0/and_13/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1617 multiplier_0/m1_n4533_n2563# multiplier_0/and_13/m1_59_58# vdd multiplier_0/and_13/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1618 multiplier_0/and_14/m1_59_58# inA1 multiplier_0/and_14/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1619 multiplier_0/and_14/nand_0/a_n5_n50# inB3 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1620 multiplier_0/and_14/m1_59_58# inA1 vdd multiplier_0/and_14/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1621 vdd inB3 multiplier_0/and_14/m1_59_58# multiplier_0/and_14/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1622 multiplier_0/m1_n4201_n2800# multiplier_0/and_14/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1623 multiplier_0/m1_n4201_n2800# multiplier_0/and_14/m1_59_58# vdd multiplier_0/and_14/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
M1624 multiplier_0/and_15/m1_59_58# inA0 multiplier_0/and_15/nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1625 multiplier_0/and_15/nand_0/a_n5_n50# inB3 gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=0 ps=0
M1626 multiplier_0/and_15/m1_59_58# inA0 vdd multiplier_0/and_15/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=0 ps=0
M1627 vdd inB3 multiplier_0/and_15/m1_59_58# multiplier_0/and_15/nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
M1628 multiplier_0/m1_n3849_n2792# multiplier_0/and_15/m1_59_58# gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=0 ps=0
M1629 multiplier_0/m1_n3849_n2792# multiplier_0/and_15/m1_59_58# vdd multiplier_0/and_15/inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=0 ps=0
C0 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# 0.63fF
C1 multiplier_0/4bitadder_0/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C2 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.13fF
C3 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_1/w_0_0# 0.04fF
C4 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n1128_n767# 0.30fF
C5 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# gnd 0.23fF
C6 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C7 vdd multiplier_0/and_10/nand_0/w_n27_n3# 0.04fF
C8 P3 gnd 0.95fF
C9 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C10 multiplier_0/4bitadder_2/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# 0.08fF
C11 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/m1_n1726_385# 0.20fF
C12 multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C13 multiplier_0/4bitadder_1/fulladder_1/m1_411_129# vdd 0.79fF
C14 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# 0.30fF
C15 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/m1_n2858_385# 0.20fF
C16 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_1/w_0_0# 0.04fF
C17 vdd multiplier_0/and_4/inverter_0/w_0_0# 0.10fF
C18 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# gnd 0.11fF
C19 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C20 gnd multiplier_0/m1_n1820_n104# 1.57fF
C21 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/m1_n2858_385# 0.08fF
C22 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C23 multiplier_0/4bitadder_0/m1_n2858_385# vdd 0.26fF
C24 multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n294_n107# 0.13fF
C25 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.30fF
C26 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# 0.13fF
C27 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/w_n27_n3# 0.13fF
C28 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# vdd 0.10fF
C29 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# gnd 0.05fF
C30 vdd multiplier_0/and_9/inverter_0/w_0_0# 0.10fF
C31 gnd multiplier_0/m1_n2968_n1347# 0.35fF
C32 inB1 multiplier_0/and_6/m1_59_58# 0.30fF
C33 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# 0.39fF
C34 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C35 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C36 vdd inA3 0.38fF
C37 vdd multiplier_0/and_13/inverter_0/w_0_0# 0.10fF
C38 gnd multiplier_0/m1_n4533_n2563# 0.46fF
C39 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n3849_n2792# 0.63fF
C40 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C41 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2617_n1342# 0.63fF
C42 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# 0.08fF
C43 multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# gnd 0.42fF
C44 multiplier_0/m1_n1473_n1361# multiplier_0/m1_n2288_n756# 1.70fF
C45 inA0 vdd 0.97fF
C46 inA3 multiplier_0/and_12/nand_0/w_n27_n3# 0.13fF
C47 inA1 inB1 1.14fF
C48 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.20fF
C49 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.13fF
C50 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C51 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# vdd 0.10fF
C52 inB2 multiplier_0/and_11/m1_59_58# 0.30fF
C53 multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# 0.03fF
C54 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n4533_n2563# 0.13fF
C55 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# 0.08fF
C56 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# 0.03fF
C57 multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# vdd 0.20fF
C58 multiplier_0/m1_n611_n78# multiplier_0/m1_n2157_n115# 3.46fF
C59 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# 0.08fF
C60 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/m1_n980_n67# 0.13fF
C61 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# 0.03fF
C62 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C63 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C64 inB0 inA2 0.86fF
C65 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# gnd 0.13fF
C66 multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# 0.20fF
C67 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C68 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_2/m1_n1726_385# 0.13fF
C69 inA1 multiplier_0/and_9/nand_0/a_n5_n50# 0.08fF
C70 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.13fF
C71 multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# 0.13fF
C72 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_0/w_0_0# 0.04fF
C73 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# 0.08fF
C74 multiplier_0/m1_n2617_n1342# multiplier_0/m1_n2968_n1347# 1.16fF
C75 multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_0/w_0_0# vdd 0.28fF
C76 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C77 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.20fF
C78 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C79 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_0/m1_n594_383# 0.13fF
C80 multiplier_0/and_4/inverter_0/w_0_0# multiplier_0/and_4/m1_59_58# 0.08fF
C81 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C82 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C83 multiplier_0/m1_n3123_n2056# gnd 2.56fF
C84 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C85 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# gnd 0.07fF
C86 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# 0.20fF
C87 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# 0.30fF
C88 multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# 0.13fF
C89 multiplier_0/m1_n3416_n801# multiplier_0/m1_n2288_n756# 6.32fF
C90 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# 0.13fF
C91 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2968_n1347# 0.63fF
C92 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n294_n107# 0.08fF
C93 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n1473_n1361# 0.30fF
C94 multiplier_0/and_14/nand_0/w_n27_n3# multiplier_0/and_14/m1_59_58# 0.13fF
C95 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# 0.20fF
C96 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# vdd 0.10fF
C97 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C98 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# 0.08fF
C99 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/a_n5_n50# 0.08fF
C100 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# 0.13fF
C101 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.13fF
C102 multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# gnd 0.09fF
C103 gnd multiplier_0/and_11/nand_0/a_n5_n50# 0.05fF
C104 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# 0.13fF
C105 multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# 0.13fF
C106 inA0 multiplier_0/and_4/m1_59_58# 0.20fF
C107 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.13fF
C108 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# 0.03fF
C109 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# 0.13fF
C110 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/m1_n594_383# 0.20fF
C111 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n2782_n115# 0.13fF
C112 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_1/w_0_0# 0.04fF
C113 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.30fF
C114 multiplier_0/and_13/inverter_0/w_0_0# multiplier_0/and_13/m1_59_58# 0.08fF
C115 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# 0.63fF
C116 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C117 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.46fF
C118 multiplier_0/m1_n2688_n2050# vdd 1.21fF
C119 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C120 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_1/m1_411_129# 0.30fF
C121 multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/w_n27_n3# vdd 0.04fF
C122 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C123 multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# vdd 0.10fF
C124 multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/w_n27_n3# vdd 0.04fF
C125 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.13fF
C126 multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# 0.03fF
C127 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C128 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C129 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# 0.03fF
C130 multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C131 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# 0.13fF
C132 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# 0.04fF
C133 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C134 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.46fF
C135 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# 0.39fF
C136 multiplier_0/4bitadder_2/m1_n594_383# gnd 0.52fF
C137 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C138 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# 0.63fF
C139 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# 0.03fF
C140 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C141 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/a_n5_n50# 0.08fF
C142 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C143 gnd multiplier_0/and_5/m1_59_58# 0.07fF
C144 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# gnd 0.05fF
C145 multiplier_0/and_6/m1_59_58# multiplier_0/m1_n2469_n98# 0.03fF
C146 multiplier_0/and_12/m1_59_58# inB3 0.30fF
C147 inB2 multiplier_0/and_10/nand_0/w_n27_n3# 0.13fF
C148 P2 gnd 3.70fF
C149 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C150 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_2/m1_411_129# 0.20fF
C151 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n980_n67# 0.13fF
C152 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# 0.20fF
C153 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_1/w_0_0# 0.04fF
C154 multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# gnd 0.09fF
C155 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C156 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# 0.03fF
C157 multiplier_0/4bitadder_1/m1_n1726_385# gnd 0.50fF
C158 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# 0.46fF
C159 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# gnd 0.07fF
C160 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# gnd 0.13fF
C161 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C162 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# vdd 0.13fF
C163 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# 0.08fF
C164 multiplier_0/m1_n294_n107# multiplier_0/m1_n1820_n104# 5.03fF
C165 inB0 multiplier_0/and_3/nand_0/w_n27_n3# 0.13fF
C166 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C167 multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# 0.08fF
C168 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# 0.63fF
C169 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_2/m1_411_129# 0.30fF
C170 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# gnd 0.05fF
C171 multiplier_0/and_15/inverter_0/w_0_0# multiplier_0/m1_n3849_n2792# 0.04fF
C172 inA3 inB2 0.83fF
C173 vdd multiplier_0/and_14/nand_0/w_n27_n3# 0.04fF
C174 vdd multiplier_0/and_3/inverter_0/w_0_0# 0.10fF
C175 gnd multiplier_0/m1_n980_n67# 7.58fF
C176 inA0 inB2 1.17fF
C177 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.13fF
C178 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# 0.13fF
C179 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n2157_n115# 0.13fF
C180 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# 0.04fF
C181 vdd multiplier_0/and_8/inverter_0/w_0_0# 0.10fF
C182 inB1 multiplier_0/and_5/m1_59_58# 0.30fF
C183 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C184 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C185 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_2/m1_n1726_385# 0.30fF
C186 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# 0.13fF
C187 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# 0.04fF
C188 multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/a_n5_n50# gnd 0.05fF
C189 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# gnd 0.26fF
C190 inA3 multiplier_0/and_7/nand_0/w_n27_n3# 0.13fF
C191 inA2 multiplier_0/and_13/nand_0/w_n27_n3# 0.13fF
C192 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# gnd 0.23fF
C193 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.13fF
C194 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.20fF
C195 multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n1820_n104# 0.30fF
C196 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# gnd 0.11fF
C197 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C198 multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C199 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n2469_n98# 0.32fF
C200 P0 vdd 7.65fF
C201 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# 0.13fF
C202 P5 gnd 1.00fF
C203 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C204 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# 0.13fF
C205 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# 0.13fF
C206 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/m1_411_129# 0.13fF
C207 multiplier_0/4bitadder_0/m1_n594_383# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# 0.08fF
C208 multiplier_0/m1_n4201_n2800# multiplier_0/m1_n3849_n2792# 1.16fF
C209 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C210 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# 0.63fF
C211 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C212 multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_1/w_0_0# gnd 0.14fF
C213 gnd multiplier_0/and_14/nand_0/a_n5_n50# 0.05fF
C214 multiplier_0/and_12/inverter_0/w_0_0# multiplier_0/and_12/m1_59_58# 0.08fF
C215 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.13fF
C216 multiplier_0/4bitadder_0/m1_n594_383# multiplier_0/4bitadder_0/halfadder_0/and_0/inverter_0/w_0_0# 0.04fF
C217 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# 0.13fF
C218 multiplier_0/and_9/nand_0/w_n27_n3# multiplier_0/and_9/m1_59_58# 0.13fF
C219 multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C220 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.20fF
C221 multiplier_0/4bitadder_1/m1_n594_383# vdd 0.36fF
C222 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.13fF
C223 multiplier_0/and_11/nand_0/w_n27_n3# multiplier_0/and_11/m1_59_58# 0.13fF
C224 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# 0.08fF
C225 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# 0.03fF
C226 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# vdd 0.79fF
C227 vdd multiplier_0/m1_n4992_n2575# 1.54fF
C228 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# 0.13fF
C229 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.30fF
C230 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C231 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C232 multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/a_n5_n50# gnd 0.05fF
C233 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n980_n67# 0.20fF
C234 inA3 multiplier_0/and_3/m1_59_58# 0.20fF
C235 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C236 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# vdd 0.10fF
C237 multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_1/w_0_0# vdd 0.13fF
C238 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# 0.04fF
C239 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n4992_n2575# 0.63fF
C240 multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# 0.63fF
C241 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.13fF
C242 multiplier_0/and_0/inverter_0/w_0_0# P0 0.04fF
C243 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/m1_n2858_385# 3.26fF
C244 multiplier_0/4bitadder_2/m1_n1726_385# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.20fF
C245 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.13fF
C246 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C247 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C248 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/m1_411_129# 0.13fF
C249 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.13fF
C250 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C251 inA0 multiplier_0/and_8/m1_59_58# 0.20fF
C252 gnd inA2 0.33fF
C253 P7 gnd 1.39fF
C254 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# 0.13fF
C255 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# 0.39fF
C256 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# gnd 0.05fF
C257 multiplier_0/4bitadder_1/m1_n2858_385# vdd 0.26fF
C258 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C259 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_1/w_0_0# 0.04fF
C260 multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n294_n107# 0.08fF
C261 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# gnd 0.13fF
C262 multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_1/w_0_0# 0.08fF
C263 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n611_n78# 0.20fF
C264 P6 gnd 1.48fF
C265 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C266 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# 0.13fF
C267 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# 0.04fF
C268 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C269 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C270 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n2157_n115# 0.32fF
C271 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C272 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C273 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/a_n5_n50# 0.08fF
C274 inB1 multiplier_0/and_4/nand_0/w_n27_n3# 0.13fF
C275 multiplier_0/and_0/m1_59_58# inA0 0.20fF
C276 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# 0.08fF
C277 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.13fF
C278 multiplier_0/and_14/inverter_0/w_0_0# multiplier_0/m1_n4201_n2800# 0.04fF
C279 vdd multiplier_0/and_12/nand_0/w_n27_n3# 0.04fF
C280 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C281 multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# vdd 0.20fF
C282 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# 0.39fF
C283 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.13fF
C284 multiplier_0/4bitadder_2/m1_n2858_385# vdd 0.26fF
C285 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C286 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C287 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C288 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/m1_n2858_385# 0.13fF
C289 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C290 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# 0.08fF
C291 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C292 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/a_n5_n50# 0.08fF
C293 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# gnd 0.05fF
C294 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.13fF
C295 multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/a_n5_n50# gnd 0.05fF
C296 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# vdd 0.04fF
C297 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C298 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C299 multiplier_0/and_10/m1_59_58# multiplier_0/m1_n3306_n1348# 0.03fF
C300 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/w_n27_n3# 0.13fF
C301 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/m1_411_129# 0.13fF
C302 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.30fF
C303 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# 0.13fF
C304 gnd multiplier_0/m1_n3602_n1349# 0.40fF
C305 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_1/w_0_0# 0.04fF
C306 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/m1_n2858_385# 0.13fF
C307 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.20fF
C308 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n3306_n1348# 0.63fF
C309 inA2 inB1 1.23fF
C310 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# vdd 0.10fF
C311 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.20fF
C312 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# 0.08fF
C313 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# 0.13fF
C314 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.13fF
C315 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/w_n27_n3# P1 0.13fF
C316 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/m1_n2858_385# 0.63fF
C317 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C318 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# 0.63fF
C319 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_0/m1_n2858_385# 0.30fF
C320 vdd multiplier_0/and_9/nand_0/w_n27_n3# 0.04fF
C321 multiplier_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C322 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_0/m1_n1726_385# 0.13fF
C323 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# 0.13fF
C324 inB2 multiplier_0/and_9/m1_59_58# 0.30fF
C325 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# 0.13fF
C326 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.20fF
C327 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/m1_n594_383# 0.20fF
C328 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C329 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C330 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_2/m1_411_129# 0.30fF
C331 multiplier_0/m1_n980_n67# multiplier_0/m1_n2469_n98# 3.46fF
C332 multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/w_n27_n3# vdd 0.04fF
C333 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/m1_n1128_n767# 0.20fF
C334 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C335 multiplier_0/and_15/m1_59_58# multiplier_0/m1_n3849_n2792# 0.03fF
C336 multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# vdd 0.10fF
C337 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/m1_n1726_385# 3.26fF
C338 inA3 multiplier_0/and_12/nand_0/a_n5_n50# 0.08fF
C339 multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# gnd 0.09fF
C340 multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/a_n5_n50# gnd 0.05fF
C341 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C342 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C343 gnd multiplier_0/m1_n2617_n1342# 0.35fF
C344 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# 0.13fF
C345 inB0 multiplier_0/and_2/m1_59_58# 0.30fF
C346 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C347 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C348 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C349 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n3602_n1349# 0.13fF
C350 multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_1/w_0_0# 0.08fF
C351 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C352 multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# gnd 0.42fF
C353 inA3 multiplier_0/and_11/nand_0/w_n27_n3# 0.13fF
C354 multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# 0.63fF
C355 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C356 gnd multiplier_0/and_4/nand_0/a_n5_n50# 0.05fF
C357 inA0 multiplier_0/and_0/nand_0/w_n27_n3# 0.13fF
C358 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C359 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.30fF
C360 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# 0.08fF
C361 multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C362 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C363 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C364 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# vdd 0.10fF
C365 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C366 multiplier_0/and_15/nand_0/w_n27_n3# multiplier_0/and_15/m1_59_58# 0.13fF
C367 gnd multiplier_0/and_9/nand_0/a_n5_n50# 0.05fF
C368 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# 0.46fF
C369 multiplier_0/4bitadder_2/m1_n594_383# multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# 0.03fF
C370 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# 0.13fF
C371 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.13fF
C372 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C373 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C374 multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/a_n5_n50# gnd 0.05fF
C375 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# 0.13fF
C376 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C377 multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_0/w_0_0# vdd 0.28fF
C378 vdd multiplier_0/m1_n611_n78# 0.90fF
C379 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/m1_n611_n78# 0.08fF
C380 multiplier_0/and_3/inverter_0/w_0_0# multiplier_0/and_3/m1_59_58# 0.08fF
C381 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C382 multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# 0.03fF
C383 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# 0.13fF
C384 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n4992_n2575# 0.13fF
C385 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_0/w_0_0# 0.04fF
C386 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/m1_n594_383# 0.13fF
C387 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/m1_n294_n107# 0.08fF
C388 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# gnd 0.27fF
C389 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# gnd 0.05fF
C390 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# gnd 0.26fF
C391 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# 0.20fF
C392 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.32fF
C393 multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_0/w_0_0# 0.08fF
C394 vdd multiplier_0/m1_n2782_n115# 1.54fF
C395 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# 0.30fF
C396 multiplier_0/and_15/nand_0/w_n27_n3# inB3 0.13fF
C397 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.13fF
C398 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# gnd 0.13fF
C399 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# gnd 0.07fF
C400 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# 0.13fF
C401 multiplier_0/m1_n4235_n2059# multiplier_0/m1_n4201_n2800# 0.24fF
C402 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# vdd 0.13fF
C403 multiplier_0/4bitadder_1/fulladder_2/m1_411_129# multiplier_0/4bitadder_1/m1_n2858_385# 3.26fF
C404 multiplier_0/and_8/inverter_0/w_0_0# multiplier_0/and_8/m1_59_58# 0.08fF
C405 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C406 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C407 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# 0.63fF
C408 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/m1_n1473_n1361# 0.20fF
C409 multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# 0.13fF
C410 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# 0.03fF
C411 multiplier_0/4bitadder_2/m1_n594_383# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.20fF
C412 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# 0.08fF
C413 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# 0.13fF
C414 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/m1_n294_n107# 0.13fF
C415 multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/m1_n1726_385# 0.13fF
C416 vdd inB2 0.81fF
C417 multiplier_0/m1_n3123_n2056# multiplier_0/m1_n3849_n2792# 10.02fF
C418 multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# 0.13fF
C419 multiplier_0/4bitadder_1/fulladder_2/m1_411_129# vdd 0.79fF
C420 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# 0.08fF
C421 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.46fF
C422 multiplier_0/4bitadder_0/fulladder_0/m1_411_129# vdd 0.79fF
C423 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.13fF
C424 gnd multiplier_0/and_12/m1_59_58# 0.07fF
C425 multiplier_0/and_11/inverter_0/w_0_0# multiplier_0/m1_n3602_n1349# 0.04fF
C426 vdd multiplier_0/and_2/nand_0/w_n27_n3# 0.04fF
C427 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C428 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# 0.08fF
C429 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.46fF
C430 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/m1_n594_383# 0.63fF
C431 multiplier_0/m1_n1473_n1361# vdd 1.39fF
C432 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# 0.04fF
C433 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/m1_n2858_385# 0.08fF
C434 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# vdd 0.13fF
C435 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# 0.03fF
C436 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C437 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_1/m1_411_129# 0.20fF
C438 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C439 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# 0.13fF
C440 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n2469_n98# 0.13fF
C441 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C442 vdd multiplier_0/and_7/nand_0/w_n27_n3# 0.04fF
C443 multiplier_0/and_5/inverter_0/w_0_0# multiplier_0/m1_n2157_n115# 0.04fF
C444 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# 0.20fF
C445 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.13fF
C446 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# 0.03fF
C447 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.30fF
C448 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C449 multiplier_0/m1_n2288_n756# multiplier_0/m1_n2968_n1347# 0.33fF
C450 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# 0.03fF
C451 vdd multiplier_0/and_1/inverter_0/w_0_0# 0.10fF
C452 multiplier_0/and_0/m1_59_58# P0 0.03fF
C453 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# 0.03fF
C454 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n3306_n1348# 0.13fF
C455 gnd multiplier_0/m1_n294_n107# 1.45fF
C456 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2782_n115# 0.63fF
C457 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/m1_n1726_385# 0.13fF
C458 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.20fF
C459 inB2 multiplier_0/and_9/nand_0/w_n27_n3# 0.13fF
C460 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# 0.13fF
C461 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# gnd 0.05fF
C462 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n1820_n104# 0.63fF
C463 multiplier_0/4bitadder_0/m1_n1726_385# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# 0.08fF
C464 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C465 multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# vdd 0.10fF
C466 vdd multiplier_0/and_6/inverter_0/w_0_0# 0.10fF
C467 gnd multiplier_0/m1_n2469_n98# 1.20fF
C468 vdd multiplier_0/and_10/inverter_0/w_0_0# 0.10fF
C469 multiplier_0/4bitadder_1/m1_n1726_385# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.20fF
C470 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C471 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# 0.13fF
C472 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C473 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.13fF
C474 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.13fF
C475 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# P1 0.30fF
C476 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C477 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/m1_n594_383# 0.20fF
C478 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# 0.08fF
C479 multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# vdd 0.20fF
C480 multiplier_0/m1_n3416_n801# vdd 1.09fF
C481 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C482 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# gnd 0.05fF
C483 multiplier_0/m1_n1128_n767# gnd 2.15fF
C484 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/m1_411_129# 0.13fF
C485 inA1 multiplier_0/and_1/nand_0/a_n5_n50# 0.08fF
C486 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_1/m1_n2858_385# 0.20fF
C487 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# 0.13fF
C488 inA3 multiplier_0/and_7/nand_0/a_n5_n50# 0.08fF
C489 multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# 0.13fF
C490 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/m1_n594_383# 3.26fF
C491 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# vdd 0.10fF
C492 multiplier_0/m1_n1820_n104# multiplier_0/m1_n2157_n115# 1.16fF
C493 multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C494 multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_1/w_0_0# vdd 0.13fF
C495 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C496 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/m1_n1726_385# 0.08fF
C497 inA2 multiplier_0/and_13/nand_0/a_n5_n50# 0.08fF
C498 multiplier_0/and_2/inverter_0/w_0_0# multiplier_0/and_2/m1_59_58# 0.08fF
C499 inA0 multiplier_0/and_0/nand_0/a_n5_n50# 0.08fF
C500 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C501 multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.20fF
C502 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# vdd 0.10fF
C503 multiplier_0/4bitadder_0/m1_n594_383# vdd 0.36fF
C504 multiplier_0/4bitadder_2/m1_n1726_385# gnd 0.50fF
C505 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# gnd 0.07fF
C506 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C507 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# 0.04fF
C508 inA1 multiplier_0/and_5/nand_0/w_n27_n3# 0.13fF
C509 multiplier_0/and_10/nand_0/w_n27_n3# multiplier_0/and_10/m1_59_58# 0.13fF
C510 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# 0.03fF
C511 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.13fF
C512 multiplier_0/m1_n2688_n2050# multiplier_0/m1_n4201_n2800# 3.46fF
C513 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C514 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# 0.13fF
C515 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_1/m1_n1726_385# 0.20fF
C516 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/a_n5_n50# 0.08fF
C517 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C518 multiplier_0/m1_n1128_n767# multiplier_0/m1_n2617_n1342# 5.03fF
C519 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n3602_n1349# 0.32fF
C520 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/a_n5_n50# 0.08fF
C521 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_0/w_0_0# 0.04fF
C522 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# 0.08fF
C523 inA2 multiplier_0/and_2/m1_59_58# 0.20fF
C524 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# 0.39fF
C525 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_0/w_0_0# 0.04fF
C526 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.13fF
C527 multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# vdd 0.20fF
C528 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# 0.08fF
C529 multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# gnd 0.09fF
C530 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C531 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C532 multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# gnd 0.09fF
C533 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C534 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/w_n27_n3# P3 0.13fF
C535 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# vdd 0.13fF
C536 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C537 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n2688_n2050# 0.13fF
C538 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/a_n5_n50# 0.08fF
C539 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C540 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C541 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_1/m1_411_129# 0.30fF
C542 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.13fF
C543 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# 0.13fF
C544 gnd multiplier_0/and_13/nand_0/a_n5_n50# 0.05fF
C545 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n3849_n2792# 0.13fF
C546 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/m1_411_129# 0.13fF
C547 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n2617_n1342# 0.13fF
C548 multiplier_0/4bitadder_1/fulladder_2/m1_411_129# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.32fF
C549 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C550 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# 0.13fF
C551 inA1 inA3 2.00fF
C552 multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_0/w_0_0# 0.08fF
C553 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.46fF
C554 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# P4 0.13fF
C555 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C556 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# 0.08fF
C557 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# gnd 0.13fF
C558 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C559 multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C560 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n4533_n2563# 0.63fF
C561 multiplier_0/and_0/m1_59_58# multiplier_0/and_0/inverter_0/w_0_0# 0.08fF
C562 multiplier_0/m1_n4235_n2059# multiplier_0/m1_n4533_n2563# 0.26fF
C563 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.46fF
C564 inA0 inA1 1.65fF
C565 inA0 multiplier_0/and_15/m1_59_58# 0.20fF
C566 multiplier_0/and_4/inverter_0/w_0_0# multiplier_0/m1_n1820_n104# 0.04fF
C567 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C568 gnd multiplier_0/and_2/m1_59_58# 0.07fF
C569 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C570 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/m1_n2858_385# 0.63fF
C571 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C572 multiplier_0/4bitadder_2/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C573 multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# vdd 0.10fF
C574 multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# 0.13fF
C575 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C576 multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.20fF
C577 inA3 inB3 0.85fF
C578 gnd multiplier_0/and_7/m1_59_58# 0.07fF
C579 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.13fF
C580 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# gnd 0.26fF
C581 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C582 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# vdd 0.10fF
C583 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C584 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# 0.13fF
C585 inA0 inB3 1.10fF
C586 multiplier_0/and_9/inverter_0/w_0_0# multiplier_0/m1_n2968_n1347# 0.04fF
C587 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.20fF
C588 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# gnd 0.13fF
C589 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n4201_n2800# 0.13fF
C590 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C591 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C592 multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_1/w_0_0# 0.08fF
C593 multiplier_0/and_13/inverter_0/w_0_0# multiplier_0/m1_n4533_n2563# 0.04fF
C594 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C595 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# gnd 0.33fF
C596 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n2968_n1347# 0.13fF
C597 multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_1/w_0_0# vdd 0.13fF
C598 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# 0.63fF
C599 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# 0.20fF
C600 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n1820_n104# 0.32fF
C601 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# 0.04fF
C602 vdd multiplier_0/and_11/nand_0/w_n27_n3# 0.04fF
C603 multiplier_0/and_5/m1_59_58# multiplier_0/m1_n2157_n115# 0.03fF
C604 vdd multiplier_0/and_0/nand_0/w_n27_n3# 0.04fF
C605 multiplier_0/m1_n4235_n2059# multiplier_0/m1_n3123_n2056# 6.32fF
C606 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C607 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# 0.13fF
C608 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/m1_411_129# 0.13fF
C609 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# 0.13fF
C610 multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# 0.03fF
C611 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C612 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C613 multiplier_0/and_14/m1_59_58# multiplier_0/m1_n4201_n2800# 0.03fF
C614 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# 0.03fF
C615 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n1473_n1361# 0.13fF
C616 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C617 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n611_n78# 0.13fF
C618 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_1/m1_411_129# 0.30fF
C619 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C620 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C621 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# gnd 0.13fF
C622 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/m1_n594_383# 0.08fF
C623 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# gnd 0.26fF
C624 multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_1/w_0_0# gnd 0.14fF
C625 multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_0/w_0_0# vdd 0.28fF
C626 gnd multiplier_0/m1_n3306_n1348# 0.38fF
C627 inB1 multiplier_0/and_7/m1_59_58# 0.30fF
C628 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# 0.04fF
C629 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.32fF
C630 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# gnd 0.05fF
C631 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C632 multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# vdd 0.10fF
C633 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# 0.13fF
C634 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.20fF
C635 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n4201_n2800# 0.30fF
C636 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C637 multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n294_n107# 0.20fF
C638 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# 0.13fF
C639 multiplier_0/4bitadder_0/m1_n1726_385# gnd 0.50fF
C640 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.13fF
C641 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.46fF
C642 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/m1_n2369_n2126# 0.13fF
C643 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# vdd 0.13fF
C644 multiplier_0/4bitadder_0/fulladder_0/m1_411_129# multiplier_0/4bitadder_0/m1_n594_383# 3.26fF
C645 vdd multiplier_0/and_15/inverter_0/w_0_0# 0.10fF
C646 gnd multiplier_0/m1_n3849_n2792# 0.46fF
C647 inB2 multiplier_0/and_8/m1_59_58# 0.30fF
C648 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/a_n5_n50# 0.08fF
C649 multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# 0.13fF
C650 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/m1_n1726_385# 0.13fF
C651 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C652 multiplier_0/m1_n980_n67# multiplier_0/m1_n2157_n115# 0.33fF
C653 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# 0.46fF
C654 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/w_n27_n3# P2 0.13fF
C655 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.30fF
C656 multiplier_0/and_5/nand_0/w_n27_n3# multiplier_0/and_5/m1_59_58# 0.13fF
C657 inB0 inA3 0.89fF
C658 multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_1/w_0_0# 0.08fF
C659 multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# vdd 0.10fF
C660 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# gnd 0.26fF
C661 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# vdd 0.04fF
C662 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C663 inA3 multiplier_0/and_11/nand_0/a_n5_n50# 0.08fF
C664 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/a_n5_n50# 0.08fF
C665 inB0 inA0 0.86fF
C666 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# 0.13fF
C667 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# 0.13fF
C668 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# 0.08fF
C669 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n2157_n115# 0.13fF
C670 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# gnd 0.26fF
C671 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C672 multiplier_0/and_1/nand_0/w_n27_n3# vdd 0.04fF
C673 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C674 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# gnd 0.05fF
C675 multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_1/w_0_0# 0.08fF
C676 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/m1_n1726_385# 0.08fF
C677 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.13fF
C678 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# 0.08fF
C679 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C680 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_0/w_0_0# 0.04fF
C681 gnd multiplier_0/and_3/nand_0/a_n5_n50# 0.05fF
C682 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C683 multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_1/w_0_0# vdd 0.13fF
C684 multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_1/w_0_0# gnd 0.14fF
C685 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# 0.08fF
C686 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/m1_n3123_n2056# 0.13fF
C687 multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C688 inA1 multiplier_0/and_14/nand_0/w_n27_n3# 0.13fF
C689 multiplier_0/and_7/inverter_0/w_0_0# multiplier_0/and_7/m1_59_58# 0.08fF
C690 vdd multiplier_0/m1_n4201_n2800# 2.94fF
C691 multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C692 gnd multiplier_0/and_8/nand_0/a_n5_n50# 0.05fF
C693 multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/m1_n1726_385# 3.26fF
C694 multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/m1_n2858_385# 0.13fF
C695 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# 0.13fF
C696 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# P3 0.30fF
C697 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/m1_n1726_385# 0.13fF
C698 multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# 0.08fF
C699 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# 0.13fF
C700 P1 vdd 5.74fF
C701 multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/w_n27_n3# vdd 0.04fF
C702 multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/a_n5_n50# gnd 0.05fF
C703 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.20fF
C704 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C705 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C706 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/m1_n2858_385# 0.20fF
C707 inA1 multiplier_0/and_9/m1_59_58# 0.20fF
C708 multiplier_0/4bitadder_1/m1_n2858_385# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.20fF
C709 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C710 multiplier_0/m1_n2688_n2050# multiplier_0/m1_n3123_n2056# 1.70fF
C711 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# 0.30fF
C712 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C713 multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_1/w_0_0# vdd 0.13fF
C714 multiplier_0/m1_n2369_n2126# gnd 2.01fF
C715 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# gnd 0.11fF
C716 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# 0.03fF
C717 multiplier_0/and_14/nand_0/w_n27_n3# inB3 0.13fF
C718 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# 0.08fF
C719 multiplier_0/4bitadder_1/fulladder_2/m1_411_129# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# 0.63fF
C720 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# 0.08fF
C721 inA1 multiplier_0/and_14/m1_59_58# 0.20fF
C722 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/m1_n2858_385# 0.08fF
C723 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C724 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.13fF
C725 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# 0.03fF
C726 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# 0.13fF
C727 multiplier_0/m1_n2288_n756# gnd 2.52fF
C728 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# 0.63fF
C729 multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2617_n1342# 0.30fF
C730 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# 0.04fF
C731 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C732 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/m1_n1726_385# 0.20fF
C733 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C734 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/m1_n594_383# 0.13fF
C735 inB2 multiplier_0/and_11/nand_0/w_n27_n3# 0.13fF
C736 multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# 0.13fF
C737 multiplier_0/4bitadder_1/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# 0.08fF
C738 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# vdd 0.10fF
C739 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_0/m1_n2858_385# 0.20fF
C740 gnd multiplier_0/and_11/m1_59_58# 0.07fF
C741 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# 0.08fF
C742 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C743 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C744 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# vdd 0.10fF
C745 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# 0.30fF
C746 multiplier_0/and_14/m1_59_58# inB3 0.30fF
C747 multiplier_0/and_9/m1_59_58# multiplier_0/m1_n2968_n1347# 0.03fF
C748 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.46fF
C749 multiplier_0/and_11/m1_59_58# multiplier_0/m1_n3602_n1349# 0.03fF
C750 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# gnd 0.07fF
C751 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C752 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# vdd 0.04fF
C753 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C754 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_0/m1_n2858_385# 0.13fF
C755 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C756 vdd multiplier_0/and_6/nand_0/w_n27_n3# 0.04fF
C757 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C758 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C759 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C760 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n4201_n2800# 0.32fF
C761 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/a_n5_n50# 0.08fF
C762 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# gnd 0.05fF
C763 multiplier_0/m1_n2288_n756# multiplier_0/m1_n2617_n1342# 10.02fF
C764 multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# 0.13fF
C765 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C766 multiplier_0/4bitadder_1/fulladder_0/m1_411_129# gnd 0.05fF
C767 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.13fF
C768 multiplier_0/4bitadder_2/m1_n2858_385# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.20fF
C769 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.46fF
C770 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/m1_n2688_n2050# 0.13fF
C771 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C772 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.20fF
C773 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# 0.08fF
C774 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# 0.13fF
C775 inA2 multiplier_0/and_6/nand_0/a_n5_n50# 0.08fF
C776 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# 0.13fF
C777 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# 0.13fF
C778 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# gnd 0.05fF
C779 multiplier_0/4bitadder_0/fulladder_0/m1_411_129# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.32fF
C780 vdd multiplier_0/and_5/inverter_0/w_0_0# 0.10fF
C781 gnd multiplier_0/m1_n2157_n115# 0.52fF
C782 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# 0.20fF
C783 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_2/m1_n1726_385# 0.20fF
C784 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/m1_n2858_385# 0.13fF
C785 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.13fF
C786 multiplier_0/and_1/inverter_0/w_0_0# multiplier_0/and_1/m1_59_58# 0.08fF
C787 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C788 P7 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# 0.20fF
C789 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# vdd 0.04fF
C790 multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# 0.08fF
C791 multiplier_0/4bitadder_0/fulladder_1/m1_411_129# gnd 0.05fF
C792 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n980_n67# 0.20fF
C793 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# 0.13fF
C794 inA0 multiplier_0/and_4/nand_0/w_n27_n3# 0.13fF
C795 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.13fF
C796 vdd inA1 0.83fF
C797 inA2 multiplier_0/and_10/nand_0/w_n27_n3# 0.13fF
C798 gnd multiplier_0/and_1/nand_0/a_n5_n50# 0.05fF
C799 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# vdd 0.10fF
C800 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C801 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# gnd 0.11fF
C802 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C803 multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/m1_n1726_385# 0.13fF
C804 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C805 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.46fF
C806 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n2369_n2126# 0.30fF
C807 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# P1 0.20fF
C808 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# 0.39fF
C809 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.13fF
C810 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C811 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C812 gnd multiplier_0/and_6/nand_0/a_n5_n50# 0.05fF
C813 inA1 multiplier_0/and_5/nand_0/a_n5_n50# 0.08fF
C814 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C815 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_1/m1_n2858_385# 0.30fF
C816 multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C817 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C818 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C819 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# 0.13fF
C820 multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_1/w_0_0# gnd 0.14fF
C821 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C822 multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# gnd 0.42fF
C823 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/m1_n2288_n756# 0.20fF
C824 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/a_n5_n50# 0.08fF
C825 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# 0.20fF
C826 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# vdd 0.10fF
C827 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C828 multiplier_0/4bitadder_1/m1_n594_383# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# 0.08fF
C829 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n2968_n1347# 0.32fF
C830 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# gnd 0.13fF
C831 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C832 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.13fF
C833 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n2157_n115# 0.13fF
C834 vdd inB3 1.01fF
C835 inA2 inA3 1.74fF
C836 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# gnd 0.26fF
C837 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C838 vdd multiplier_0/m1_n1820_n104# 1.31fF
C839 multiplier_0/m1_n4235_n2059# gnd 2.47fF
C840 inA0 inA2 1.66fF
C841 multiplier_0/and_12/nand_0/w_n27_n3# inB3 0.13fF
C842 inA1 multiplier_0/and_9/nand_0/w_n27_n3# 0.13fF
C843 multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/a_n5_n50# gnd 0.05fF
C844 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C845 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C846 vdd multiplier_0/m1_n2968_n1347# 2.94fF
C847 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# 0.13fF
C848 multiplier_0/and_0/m1_59_58# multiplier_0/and_0/nand_0/w_n27_n3# 0.13fF
C849 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# vdd 0.10fF
C850 vdd multiplier_0/m1_n4533_n2563# 1.54fF
C851 multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_0/w_0_0# vdd 0.28fF
C852 multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# vdd 0.10fF
C853 multiplier_0/4bitadder_1/fulladder_1/m1_411_129# gnd 0.05fF
C854 multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_0/w_0_0# 0.08fF
C855 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.46fF
C856 multiplier_0/4bitadder_1/fulladder_0/m1_411_129# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.32fF
C857 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C858 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C859 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C860 multiplier_0/4bitadder_0/m1_n2858_385# gnd 0.50fF
C861 multiplier_0/and_11/inverter_0/w_0_0# multiplier_0/and_11/m1_59_58# 0.08fF
C862 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# 0.13fF
C863 multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# 0.20fF
C864 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# 0.20fF
C865 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# gnd 0.07fF
C866 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C867 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n3602_n1349# 0.63fF
C868 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C869 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_1/m1_411_129# 0.20fF
C870 gnd inA3 0.33fF
C871 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C872 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C873 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n611_n78# 0.20fF
C874 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_0/m1_411_129# 0.30fF
C875 multiplier_0/and_3/inverter_0/w_0_0# multiplier_0/m1_n980_n67# 0.04fF
C876 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# P4 0.30fF
C877 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# 0.08fF
C878 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/m1_411_129# 0.13fF
C879 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# gnd 0.26fF
C880 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/m1_n594_383# 0.13fF
C881 multiplier_0/and_12/inverter_0/w_0_0# multiplier_0/m1_n4992_n2575# 0.04fF
C882 inA0 gnd 0.33fF
C883 inB1 multiplier_0/and_5/nand_0/w_n27_n3# 0.13fF
C884 multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# gnd 0.09fF
C885 multiplier_0/and_4/m1_59_58# multiplier_0/m1_n1820_n104# 0.03fF
C886 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_1/m1_411_129# 0.30fF
C887 multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n3849_n2792# 0.30fF
C888 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C889 multiplier_0/m1_n3123_n2056# vdd 1.21fF
C890 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n294_n107# 0.63fF
C891 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C892 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n611_n78# 0.08fF
C893 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C894 multiplier_0/4bitadder_0/m1_n2858_385# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# 0.08fF
C895 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# 0.04fF
C896 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C897 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# 0.20fF
C898 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# 0.13fF
C899 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n2469_n98# 0.13fF
C900 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# 0.13fF
C901 inB0 vdd 1.37fF
C902 multiplier_0/and_13/m1_59_58# inB3 0.30fF
C903 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# 0.13fF
C904 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# gnd 0.23fF
C905 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# 0.20fF
C906 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.46fF
C907 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# P6 0.13fF
C908 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# 0.08fF
C909 multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# vdd 0.20fF
C910 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# 0.03fF
C911 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# 0.13fF
C912 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# 0.04fF
C913 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# 0.20fF
C914 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/m1_n1726_385# 0.08fF
C915 vdd multiplier_0/and_12/inverter_0/w_0_0# 0.10fF
C916 P4 gnd 0.90fF
C917 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.13fF
C918 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# multiplier_0/m1_n980_n67# 0.08fF
C919 multiplier_0/and_13/m1_59_58# multiplier_0/m1_n4533_n2563# 0.03fF
C920 inA3 inB1 1.02fF
C921 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/m1_n2858_385# 0.08fF
C922 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.13fF
C923 inB2 multiplier_0/and_10/m1_59_58# 0.30fF
C924 inA0 inB1 1.34fF
C925 multiplier_0/4bitadder_2/m1_n1726_385# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# 0.08fF
C926 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.30fF
C927 multiplier_0/m1_n611_n78# multiplier_0/m1_n1820_n104# 0.28fF
C928 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_0/w_0_0# 0.04fF
C929 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C930 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.13fF
C931 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# 0.08fF
C932 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# vdd 0.04fF
C933 inA1 inB2 1.18fF
C934 inA0 multiplier_0/and_4/nand_0/a_n5_n50# 0.08fF
C935 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# 0.08fF
C936 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# 0.13fF
C937 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# 0.13fF
C938 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/m1_n1726_385# 0.13fF
C939 inA2 multiplier_0/and_10/nand_0/a_n5_n50# 0.08fF
C940 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C941 multiplier_0/4bitadder_2/m1_n594_383# vdd 0.36fF
C942 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n4201_n2800# 0.63fF
C943 multiplier_0/4bitadder_1/fulladder_2/m1_411_129# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C944 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C945 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# vdd 0.79fF
C946 multiplier_0/m1_n2688_n2050# gnd 2.01fF
C947 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C948 multiplier_0/and_3/nand_0/w_n27_n3# inA3 0.13fF
C949 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_2/m1_n594_383# 0.13fF
C950 P2 vdd 3.25fF
C951 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C952 multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# gnd 0.42fF
C953 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C954 multiplier_0/4bitadder_0/m1_n2858_385# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.20fF
C955 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/m1_411_129# 0.63fF
C956 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C957 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# 0.13fF
C958 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/w_n27_n3# 0.13fF
C959 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# 0.13fF
C960 multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/w_n27_n3# vdd 0.04fF
C961 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# gnd 0.23fF
C962 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C963 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# P5 0.13fF
C964 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# 0.08fF
C965 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# 0.13fF
C966 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# 0.03fF
C967 inA0 multiplier_0/and_8/nand_0/w_n27_n3# 0.13fF
C968 multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# vdd 0.20fF
C969 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n2782_n115# 0.13fF
C970 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# 0.20fF
C971 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.13fF
C972 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/m1_n1726_385# 0.08fF
C973 multiplier_0/4bitadder_1/m1_n1726_385# vdd 0.26fF
C974 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/m1_n2369_n2126# 0.20fF
C975 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# P2 0.30fF
C976 multiplier_0/and_6/inverter_0/w_0_0# multiplier_0/and_6/m1_59_58# 0.08fF
C977 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# 0.63fF
C978 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# 0.13fF
C979 multiplier_0/and_10/inverter_0/w_0_0# multiplier_0/and_10/m1_59_58# 0.08fF
C980 gnd multiplier_0/and_10/nand_0/a_n5_n50# 0.05fF
C981 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/m1_n2858_385# 0.08fF
C982 multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_0/w_0_0# vdd 0.28fF
C983 vdd multiplier_0/m1_n980_n67# 0.84fF
C984 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# 0.08fF
C985 multiplier_0/m1_n1473_n1361# multiplier_0/m1_n2968_n1347# 3.46fF
C986 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C987 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# vdd 0.04fF
C988 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.13fF
C989 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# gnd 0.07fF
C990 gnd multiplier_0/and_15/nand_0/a_n5_n50# 0.05fF
C991 inA3 multiplier_0/and_12/m1_59_58# 0.20fF
C992 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C993 multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.32fF
C994 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# gnd 0.05fF
C995 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C996 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.13fF
C997 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# 0.13fF
C998 multiplier_0/and_1/nand_0/w_n27_n3# multiplier_0/and_1/m1_59_58# 0.13fF
C999 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C1000 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/m1_n2858_385# 0.13fF
C1001 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C1002 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C1003 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# vdd 0.10fF
C1004 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1005 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C1006 multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_1/w_0_0# 0.08fF
C1007 multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_0/w_0_0# 0.08fF
C1008 multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# 0.13fF
C1009 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C1010 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# 0.13fF
C1011 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n3123_n2056# 0.30fF
C1012 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/m1_n2858_385# 0.13fF
C1013 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C1014 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1015 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# vdd 0.10fF
C1016 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1017 gnd multiplier_0/and_9/m1_59_58# 0.07fF
C1018 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# P3 0.20fF
C1019 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/m1_n2858_385# 0.63fF
C1020 multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/w_n27_n3# vdd 0.04fF
C1021 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n2968_n1347# 0.13fF
C1022 multiplier_0/4bitadder_0/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# 0.08fF
C1023 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# 0.08fF
C1024 multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# 0.13fF
C1025 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/m1_n2858_385# 3.26fF
C1026 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n4992_n2575# 0.30fF
C1027 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_2/m1_n2858_385# 0.30fF
C1028 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_1/w_0_0# 0.04fF
C1029 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.30fF
C1030 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# vdd 0.04fF
C1031 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C1032 multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_1/w_0_0# vdd 0.13fF
C1033 vdd multiplier_0/and_4/nand_0/w_n27_n3# 0.04fF
C1034 multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C1035 multiplier_0/m1_n3416_n801# multiplier_0/m1_n2968_n1347# 0.24fF
C1036 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1037 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/m1_n594_383# 0.63fF
C1038 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C1039 gnd multiplier_0/and_14/m1_59_58# 0.07fF
C1040 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C1041 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C1042 inB0 multiplier_0/and_2/nand_0/w_n27_n3# 0.13fF
C1043 P0 gnd 7.92fF
C1044 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.46fF
C1045 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C1046 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# 0.39fF
C1047 multiplier_0/m1_n2288_n756# multiplier_0/m1_n3306_n1348# 3.46fF
C1048 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C1049 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/a_n5_n50# 0.08fF
C1050 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/m1_n611_n78# 0.13fF
C1051 vdd multiplier_0/and_13/nand_0/w_n27_n3# 0.04fF
C1052 vdd multiplier_0/and_2/inverter_0/w_0_0# 0.10fF
C1053 multiplier_0/m1_n2369_n2126# multiplier_0/m1_n3849_n2792# 5.03fF
C1054 multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_1/w_0_0# 0.08fF
C1055 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C1056 multiplier_0/and_8/inverter_0/w_0_0# multiplier_0/m1_n2617_n1342# 0.04fF
C1057 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/w_n27_n3# 0.13fF
C1058 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/m1_n594_383# 0.08fF
C1059 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/m1_n594_383# 0.08fF
C1060 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n4533_n2563# 0.13fF
C1061 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1062 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C1063 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.20fF
C1064 multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# 0.03fF
C1065 multiplier_0/4bitadder_1/m1_n594_383# gnd 0.52fF
C1066 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C1067 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# 0.13fF
C1068 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1069 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C1070 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C1071 vdd inA2 0.86fF
C1072 gnd multiplier_0/m1_n4992_n2575# 0.54fF
C1073 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# gnd 0.05fF
C1074 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# vdd 0.13fF
C1075 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1076 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C1077 multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n2617_n1342# 0.13fF
C1078 multiplier_0/m1_n611_n78# multiplier_0/m1_n980_n67# 1.70fF
C1079 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C1080 multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_1/w_0_0# gnd 0.14fF
C1081 multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_0/w_0_0# vdd 0.28fF
C1082 multiplier_0/4bitadder_2/m1_n594_383# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# 0.08fF
C1083 multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# 0.08fF
C1084 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2469_n98# 0.30fF
C1085 multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_0/w_0_0# 0.08fF
C1086 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.46fF
C1087 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/m1_n2288_n756# 0.13fF
C1088 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C1089 multiplier_0/4bitadder_0/fulladder_1/m1_411_129# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C1090 multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# 0.04fF
C1091 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.46fF
C1092 multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n3849_n2792# 0.13fF
C1093 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1094 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n2688_n2050# 0.30fF
C1095 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# gnd 0.07fF
C1096 multiplier_0/and_4/nand_0/w_n27_n3# multiplier_0/and_4/m1_59_58# 0.13fF
C1097 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# 0.13fF
C1098 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# 0.13fF
C1099 multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# 0.13fF
C1100 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C1101 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C1102 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# gnd 0.13fF
C1103 multiplier_0/4bitadder_1/m1_n2858_385# gnd 0.50fF
C1104 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.13fF
C1105 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/m1_n1726_385# 0.63fF
C1106 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C1107 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C1108 P7 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# 0.30fF
C1109 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# gnd 0.05fF
C1110 inB0 multiplier_0/and_3/m1_59_58# 0.30fF
C1111 multiplier_0/4bitadder_1/m1_n594_383# multiplier_0/4bitadder_1/halfadder_0/and_0/inverter_0/w_0_0# 0.04fF
C1112 gnd vdd 10.13fF
C1113 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C1114 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# 0.13fF
C1115 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.46fF
C1116 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n4201_n2800# 0.13fF
C1117 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C1118 multiplier_0/4bitadder_0/fulladder_1/m1_411_129# multiplier_0/4bitadder_0/m1_n1726_385# 3.26fF
C1119 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C1120 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/m1_n594_383# 0.08fF
C1121 vdd multiplier_0/m1_n3602_n1349# 1.54fF
C1122 multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# gnd 0.09fF
C1123 gnd multiplier_0/and_5/nand_0/a_n5_n50# 0.05fF
C1124 multiplier_0/4bitadder_2/m1_n2858_385# gnd 0.50fF
C1125 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C1126 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n4533_n2563# 0.13fF
C1127 multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_0/w_0_0# multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# 0.08fF
C1128 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1129 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# gnd 0.13fF
C1130 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2157_n115# 0.63fF
C1131 multiplier_0/and_13/nand_0/w_n27_n3# multiplier_0/and_13/m1_59_58# 0.13fF
C1132 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/w_n27_n3# 0.13fF
C1133 inA1 multiplier_0/and_1/m1_59_58# 0.20fF
C1134 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C1135 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_1/w_0_0# 0.04fF
C1136 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# 0.13fF
C1137 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C1138 multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/a_n5_n50# gnd 0.05fF
C1139 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# 0.20fF
C1140 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.20fF
C1141 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# 0.08fF
C1142 inA3 multiplier_0/and_7/m1_59_58# 0.20fF
C1143 inB0 multiplier_0/and_0/m1_59_58# 0.30fF
C1144 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/m1_411_129# 0.13fF
C1145 multiplier_0/4bitadder_1/m1_n1726_385# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# 0.08fF
C1146 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# 0.30fF
C1147 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# 0.39fF
C1148 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# 0.08fF
C1149 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# 0.03fF
C1150 inA2 multiplier_0/and_13/m1_59_58# 0.20fF
C1151 multiplier_0/and_2/inverter_0/w_0_0# multiplier_0/m1_n611_n78# 0.04fF
C1152 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# gnd 0.11fF
C1153 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# 0.04fF
C1154 multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# vdd 0.20fF
C1155 vdd multiplier_0/m1_n2617_n1342# 1.31fF
C1156 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C1157 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n3306_n1348# 0.13fF
C1158 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/a_n5_n50# 0.08fF
C1159 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n1820_n104# 0.13fF
C1160 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_0/w_0_0# 0.04fF
C1161 multiplier_0/and_15/inverter_0/w_0_0# multiplier_0/and_15/m1_59_58# 0.08fF
C1162 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.20fF
C1163 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# vdd 0.10fF
C1164 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# 0.03fF
C1165 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_1/m1_n1726_385# 0.13fF
C1166 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# 0.20fF
C1167 multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# vdd 0.10fF
C1168 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C1169 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/w_n27_n3# 0.13fF
C1170 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/m1_411_129# 0.13fF
C1171 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.32fF
C1172 vdd inB1 2.47fF
C1173 multiplier_0/m1_n4235_n2059# multiplier_0/m1_n3849_n2792# 0.22fF
C1174 multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# gnd 0.42fF
C1175 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n2617_n1342# 0.13fF
C1176 multiplier_0/4bitadder_1/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C1177 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_0/w_0_0# 0.04fF
C1178 gnd multiplier_0/and_4/m1_59_58# 0.07fF
C1179 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# 0.13fF
C1180 multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# 0.08fF
C1181 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C1182 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n2617_n1342# 0.32fF
C1183 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# 0.13fF
C1184 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# gnd 0.86fF
C1185 multiplier_0/4bitadder_0/fulladder_0/m1_411_129# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C1186 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.20fF
C1187 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C1188 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# 0.20fF
C1189 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C1190 multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/m1_n2858_385# 0.13fF
C1191 multiplier_0/4bitadder_0/m1_n594_383# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.20fF
C1192 multiplier_0/and_1/nand_0/w_n27_n3# inA1 0.13fF
C1193 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1194 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C1195 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C1196 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n2782_n115# 0.13fF
C1197 multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_1/w_0_0# 0.08fF
C1198 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# 0.13fF
C1199 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n2782_n115# 0.32fF
C1200 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n980_n67# 0.08fF
C1201 gnd multiplier_0/and_13/m1_59_58# 0.07fF
C1202 vdd multiplier_0/and_3/nand_0/w_n27_n3# 0.04fF
C1203 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C1204 multiplier_0/and_3/m1_59_58# multiplier_0/m1_n980_n67# 0.03fF
C1205 multiplier_0/and_12/m1_59_58# multiplier_0/m1_n4992_n2575# 0.03fF
C1206 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.13fF
C1207 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.32fF
C1208 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# P4 0.20fF
C1209 multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/w_n27_n3# vdd 0.04fF
C1210 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# 0.08fF
C1211 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# gnd 0.11fF
C1212 vdd multiplier_0/and_8/nand_0/w_n27_n3# 0.04fF
C1213 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# vdd 0.13fF
C1214 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C1215 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# vdd 0.10fF
C1216 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# 0.03fF
C1217 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_0/m1_n1726_385# 0.20fF
C1218 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C1219 inA2 inB2 1.02fF
C1220 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1221 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/m1_n1726_385# 0.63fF
C1222 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/w_n27_n3# 0.13fF
C1223 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.13fF
C1224 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C1225 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# 0.03fF
C1226 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C1227 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C1228 gnd multiplier_0/m1_n611_n78# 1.45fF
C1229 multiplier_0/and_2/nand_0/w_n27_n3# inA2 0.13fF
C1230 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.30fF
C1231 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n2968_n1347# 0.13fF
C1232 vdd multiplier_0/and_7/inverter_0/w_0_0# 0.10fF
C1233 inB1 multiplier_0/and_4/m1_59_58# 0.30fF
C1234 inB0 multiplier_0/and_0/nand_0/w_n27_n3# 0.13fF
C1235 multiplier_0/4bitadder_2/m1_n594_383# multiplier_0/4bitadder_2/halfadder_0/and_0/inverter_0/w_0_0# 0.04fF
C1236 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1237 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# 0.13fF
C1238 gnd multiplier_0/m1_n2782_n115# 4.24fF
C1239 vdd multiplier_0/and_11/inverter_0/w_0_0# 0.10fF
C1240 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# P6 0.30fF
C1241 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C1242 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/m1_411_129# 0.13fF
C1243 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n980_n67# 0.13fF
C1244 inB0 multiplier_0/and_1/m1_59_58# 0.30fF
C1245 multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n1820_n104# 0.13fF
C1246 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# gnd 0.05fF
C1247 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# 0.13fF
C1248 inA3 multiplier_0/and_3/nand_0/a_n5_n50# 0.08fF
C1249 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# 0.13fF
C1250 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/m1_n1726_385# 0.13fF
C1251 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C1252 multiplier_0/and_12/nand_0/w_n27_n3# multiplier_0/and_12/m1_59_58# 0.13fF
C1253 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_1/m1_n2858_385# 0.13fF
C1254 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.13fF
C1255 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# 0.08fF
C1256 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.13fF
C1257 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# vdd 0.04fF
C1258 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n4533_n2563# 0.30fF
C1259 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# 0.04fF
C1260 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/m1_n1726_385# 0.08fF
C1261 multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# 0.08fF
C1262 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/m1_n2858_385# 0.13fF
C1263 multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# 0.13fF
C1264 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C1265 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C1266 multiplier_0/4bitadder_1/fulladder_2/m1_411_129# gnd 0.05fF
C1267 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/m1_n2688_n2050# 0.20fF
C1268 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n980_n67# 0.63fF
C1269 multiplier_0/4bitadder_0/fulladder_0/m1_411_129# gnd 0.05fF
C1270 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/m1_n594_383# 0.13fF
C1271 inA0 multiplier_0/and_15/nand_0/w_n27_n3# 0.13fF
C1272 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1273 multiplier_0/m1_n1473_n1361# gnd 2.20fF
C1274 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C1275 multiplier_0/4bitadder_0/fulladder_1/m1_411_129# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.32fF
C1276 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n611_n78# 0.13fF
C1277 inA0 multiplier_0/and_8/nand_0/a_n5_n50# 0.08fF
C1278 multiplier_0/and_6/nand_0/w_n27_n3# multiplier_0/and_6/m1_59_58# 0.13fF
C1279 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C1280 vdd multiplier_0/m1_n294_n107# 0.61fF
C1281 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# gnd 0.05fF
C1282 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# 0.03fF
C1283 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# vdd 0.13fF
C1284 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C1285 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.13fF
C1286 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C1287 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# 0.03fF
C1288 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2968_n1347# 0.30fF
C1289 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# vdd 0.10fF
C1290 multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C1291 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# 0.08fF
C1292 vdd multiplier_0/m1_n2469_n98# 1.54fF
C1293 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/a_n5_n50# 0.08fF
C1294 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.13fF
C1295 multiplier_0/m1_n2688_n2050# multiplier_0/m1_n3849_n2792# 0.28fF
C1296 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_1/m1_411_129# 0.30fF
C1297 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C1298 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# P5 0.30fF
C1299 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# 0.13fF
C1300 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.13fF
C1301 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/m1_n1726_385# 0.63fF
C1302 multiplier_0/and_1/nand_0/w_n27_n3# inB0 0.13fF
C1303 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1304 multiplier_0/m1_n1128_n767# vdd 1.14fF
C1305 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C1306 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# 0.03fF
C1307 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# vdd 0.79fF
C1308 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C1309 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n4533_n2563# 0.32fF
C1310 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# P2 0.20fF
C1311 multiplier_0/m1_n3123_n2056# multiplier_0/m1_n4201_n2800# 0.33fF
C1312 multiplier_0/m1_n3123_n2056# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# 0.20fF
C1313 multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# gnd 0.42fF
C1314 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C1315 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# 0.39fF
C1316 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_2/m1_n2858_385# 0.13fF
C1317 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C1318 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# gnd 0.05fF
C1319 multiplier_0/m1_n1473_n1361# multiplier_0/m1_n2617_n1342# 0.28fF
C1320 inA3 multiplier_0/and_11/m1_59_58# 0.20fF
C1321 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/w_n27_n3# 0.13fF
C1322 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2782_n115# 0.30fF
C1323 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# 0.13fF
C1324 multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# gnd 0.09fF
C1325 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# 0.08fF
C1326 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# 0.13fF
C1327 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1328 multiplier_0/4bitadder_1/m1_n594_383# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.20fF
C1329 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# gnd 0.23fF
C1330 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# 0.13fF
C1331 multiplier_0/m1_n3416_n801# gnd 2.32fF
C1332 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# 0.13fF
C1333 multiplier_0/4bitadder_2/m1_n1726_385# vdd 0.26fF
C1334 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# 0.13fF
C1335 multiplier_0/m1_n3416_n801# multiplier_0/m1_n3602_n1349# 3.96fF
C1336 multiplier_0/m1_n1473_n1361# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# 0.63fF
C1337 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.30fF
C1338 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C1339 multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_0/w_0_0# 0.08fF
C1340 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.46fF
C1341 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/m1_n1128_n767# 0.13fF
C1342 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# 0.13fF
C1343 inB1 multiplier_0/and_7/nand_0/w_n27_n3# 0.13fF
C1344 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C1345 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# 0.30fF
C1346 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# vdd 0.13fF
C1347 multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_1/w_0_0# gnd 0.14fF
C1348 multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_0/w_0_0# vdd 0.28fF
C1349 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# 0.20fF
C1350 gnd multiplier_0/and_3/m1_59_58# 0.07fF
C1351 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n3849_n2792# 0.13fF
C1352 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.30fF
C1353 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# 0.13fF
C1354 inB2 multiplier_0/and_8/nand_0/w_n27_n3# 0.13fF
C1355 multiplier_0/and_7/inverter_0/w_0_0# multiplier_0/m1_n2782_n115# 0.04fF
C1356 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n3849_n2792# 0.32fF
C1357 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/m1_n3123_n2056# 0.20fF
C1358 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# gnd 0.26fF
C1359 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/m1_n594_383# 0.08fF
C1360 multiplier_0/4bitadder_0/m1_n594_383# gnd 0.52fF
C1361 gnd multiplier_0/and_8/m1_59_58# 0.07fF
C1362 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C1363 multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# vdd 0.20fF
C1364 multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# vdd 0.20fF
C1365 inA1 inB3 1.24fF
C1366 inB3 multiplier_0/and_15/m1_59_58# 0.30fF
C1367 multiplier_0/and_0/m1_59_58# gnd 0.07fF
C1368 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C1369 multiplier_0/m1_n3416_n801# multiplier_0/m1_n2617_n1342# 0.22fF
C1370 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C1371 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# vdd 0.10fF
C1372 multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# 0.13fF
C1373 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.13fF
C1374 multiplier_0/m1_n294_n107# multiplier_0/m1_n611_n78# 0.59fF
C1375 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# gnd 0.23fF
C1376 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/m1_n294_n107# 0.20fF
C1377 multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# gnd 0.09fF
C1378 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C1379 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# 0.13fF
C1380 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# multiplier_0/m1_n980_n67# 0.08fF
C1381 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# gnd 0.05fF
C1382 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# 0.03fF
C1383 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n3602_n1349# 0.13fF
C1384 multiplier_0/and_8/m1_59_58# multiplier_0/m1_n2617_n1342# 0.03fF
C1385 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_2/m1_n1726_385# 0.08fF
C1386 multiplier_0/4bitadder_1/m1_n2858_385# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# 0.08fF
C1387 multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# 0.03fF
C1388 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# 0.08fF
C1389 multiplier_0/m1_n4235_n2059# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# 0.13fF
C1390 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.30fF
C1391 multiplier_0/4bitadder_1/fulladder_1/m1_411_129# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C1392 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C1393 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C1394 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# 0.30fF
C1395 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# vdd 0.10fF
C1396 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# 0.13fF
C1397 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# multiplier_0/4bitadder_0/m1_n594_383# 0.08fF
C1398 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# 0.13fF
C1399 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# 0.08fF
C1400 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C1401 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/m1_n594_383# 0.13fF
C1402 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# gnd 0.05fF
C1403 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1404 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.20fF
C1405 multiplier_0/m1_n3416_n801# multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# 0.20fF
C1406 multiplier_0/and_3/nand_0/w_n27_n3# multiplier_0/and_3/m1_59_58# 0.13fF
C1407 multiplier_0/m1_n2369_n2126# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C1408 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n3306_n1348# 0.13fF
C1409 multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# gnd 0.42fF
C1410 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n4992_n2575# 0.13fF
C1411 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.13fF
C1412 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/m1_n1473_n1361# 0.13fF
C1413 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C1414 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_1/w_0_0# 0.04fF
C1415 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# multiplier_0/m1_n2288_n756# 0.30fF
C1416 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# gnd 0.23fF
C1417 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.13fF
C1418 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.05fF
C1419 multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/w_n27_n3# vdd 0.04fF
C1420 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# gnd 0.23fF
C1421 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# gnd 0.11fF
C1422 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C1423 multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# 0.13fF
C1424 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# 0.08fF
C1425 inB0 inA1 0.85fF
C1426 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/m1_n594_383# 0.63fF
C1427 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# 0.08fF
C1428 multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# 0.13fF
C1429 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# multiplier_0/4bitadder_1/m1_n2858_385# 0.08fF
C1430 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_1/m1_n1726_385# 0.30fF
C1431 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.20fF
C1432 gnd multiplier_0/and_12/nand_0/a_n5_n50# 0.05fF
C1433 multiplier_0/and_8/nand_0/w_n27_n3# multiplier_0/and_8/m1_59_58# 0.13fF
C1434 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.13fF
C1435 multiplier_0/and_1/inverter_0/w_0_0# multiplier_0/m1_n294_n107# 0.04fF
C1436 multiplier_0/4bitadder_0/m1_n1726_385# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.20fF
C1437 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# 0.08fF
C1438 inA0 inA3 1.72fF
C1439 multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_1/w_0_0# gnd 0.14fF
C1440 multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_0/w_0_0# vdd 0.28fF
C1441 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# vdd 0.10fF
C1442 multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_1/w_0_0# vdd 0.13fF
C1443 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_1/m1_n1726_385# 0.13fF
C1444 multiplier_0/4bitadder_0/fulladder_1/m1_411_129# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# 0.63fF
C1445 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.13fF
C1446 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C1447 multiplier_0/and_5/inverter_0/w_0_0# multiplier_0/and_5/m1_59_58# 0.08fF
C1448 multiplier_0/4bitadder_2/m1_n2858_385# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# 0.08fF
C1449 vdd multiplier_0/m1_n3306_n1348# 1.54fF
C1450 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.13fF
C1451 multiplier_0/and_14/inverter_0/w_0_0# multiplier_0/and_14/m1_59_58# 0.08fF
C1452 gnd multiplier_0/and_1/m1_59_58# 0.07fF
C1453 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1454 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# multiplier_0/4bitadder_2/m1_n2858_385# 0.20fF
C1455 multiplier_0/4bitadder_1/m1_n594_383# multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# 0.03fF
C1456 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C1457 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# 0.30fF
C1458 multiplier_0/4bitadder_0/m1_n1726_385# vdd 0.26fF
C1459 vdd multiplier_0/m1_n3849_n2792# 1.31fF
C1460 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# gnd 0.07fF
C1461 multiplier_0/m1_n3123_n2056# multiplier_0/m1_n4533_n2563# 3.46fF
C1462 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# 0.03fF
C1463 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# 0.08fF
C1464 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# 0.13fF
C1465 multiplier_0/and_6/inverter_0/w_0_0# multiplier_0/m1_n2469_n98# 0.04fF
C1466 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# 0.13fF
C1467 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C1468 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# 0.30fF
C1469 inA1 multiplier_0/and_5/m1_59_58# 0.20fF
C1470 multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_1/w_0_0# 0.08fF
C1471 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# 0.13fF
C1472 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C1473 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_2/m1_411_129# 0.30fF
C1474 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# 0.30fF
C1475 multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# gnd 0.42fF
C1476 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# vdd 0.10fF
C1477 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_0/w_0_0# 0.04fF
C1478 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n4201_n2800# 0.13fF
C1479 multiplier_0/and_2/m1_59_58# multiplier_0/m1_n611_n78# 0.03fF
C1480 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C1481 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C1482 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# vdd 0.10fF
C1483 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C1484 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# gnd 0.05fF
C1485 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n2157_n115# 0.30fF
C1486 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# vdd 0.79fF
C1487 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C1488 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# 0.03fF
C1489 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.13fF
C1490 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.30fF
C1491 multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# gnd 0.42fF
C1492 multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_1/w_0_0# vdd 0.13fF
C1493 multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_0/w_0_0# 0.08fF
C1494 multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_0/m1_n1726_385# 0.13fF
C1495 vdd multiplier_0/and_15/nand_0/w_n27_n3# 0.04fF
C1496 multiplier_0/and_7/m1_59_58# multiplier_0/m1_n2782_n115# 0.03fF
C1497 P7 multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/w_n27_n3# 0.13fF
C1498 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C1499 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# 0.13fF
C1500 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_1/m1_n594_383# 0.13fF
C1501 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1502 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.30fF
C1503 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C1504 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C1505 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n3306_n1348# 0.30fF
C1506 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C1507 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# 0.30fF
C1508 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# 0.20fF
C1509 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# vdd 0.04fF
C1510 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C1511 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C1512 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C1513 multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_1/w_0_0# gnd 0.14fF
C1514 multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_0/w_0_0# vdd 0.28fF
C1515 vdd multiplier_0/and_14/inverter_0/w_0_0# 0.10fF
C1516 gnd multiplier_0/m1_n4201_n2800# 0.46fF
C1517 inA2 multiplier_0/and_2/nand_0/a_n5_n50# 0.08fF
C1518 multiplier_0/and_2/nand_0/w_n27_n3# multiplier_0/and_2/m1_59_58# 0.13fF
C1519 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_2/m1_411_129# 0.30fF
C1520 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C1521 multiplier_0/4bitadder_1/fulladder_0/m1_411_129# multiplier_0/4bitadder_1/m1_n594_383# 3.26fF
C1522 multiplier_0/4bitadder_0/m1_n594_383# multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# 0.03fF
C1523 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n2469_n98# 0.13fF
C1524 multiplier_0/m1_n2369_n2126# vdd 1.00fF
C1525 multiplier_0/m1_n980_n67# multiplier_0/m1_n1820_n104# 10.02fF
C1526 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# vdd 0.10fF
C1527 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C1528 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# multiplier_0/4bitadder_0/m1_n1726_385# 0.30fF
C1529 multiplier_0/m1_n2288_n756# vdd 1.19fF
C1530 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# gnd 0.05fF
C1531 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# 0.08fF
C1532 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# 0.13fF
C1533 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C1534 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# 0.04fF
C1535 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C1536 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n3306_n1348# 0.32fF
C1537 P1 gnd 6.36fF
C1538 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C1539 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C1540 multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# 0.13fF
C1541 multiplier_0/and_7/nand_0/w_n27_n3# multiplier_0/and_7/m1_59_58# 0.13fF
C1542 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# gnd 0.05fF
C1543 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.13fF
C1544 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C1545 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# gnd 0.13fF
C1546 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n2469_n98# 0.63fF
C1547 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# gnd 0.05fF
C1548 inA2 multiplier_0/and_6/nand_0/w_n27_n3# 0.13fF
C1549 multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/w_n27_n3# vdd 0.04fF
C1550 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# 0.30fF
C1551 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# gnd 0.07fF
C1552 multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_1/w_0_0# gnd 0.14fF
C1553 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1554 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1555 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.13fF
C1556 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# P6 0.20fF
C1557 inA1 multiplier_0/and_14/nand_0/a_n5_n50# 0.08fF
C1558 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# 0.13fF
C1559 inA0 multiplier_0/and_15/nand_0/a_n5_n50# 0.08fF
C1560 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# multiplier_0/m1_n3602_n1349# 0.30fF
C1561 gnd multiplier_0/and_2/nand_0/a_n5_n50# 0.05fF
C1562 multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/m1_n2858_385# 0.13fF
C1563 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# 0.20fF
C1564 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# 0.13fF
C1565 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# gnd 0.13fF
C1566 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# 0.30fF
C1567 multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# 0.04fF
C1568 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# multiplier_0/4bitadder_1/fulladder_0/m1_411_129# 0.30fF
C1569 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C1570 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C1571 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/m1_n611_n78# 0.63fF
C1572 multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/w_n27_n3# vdd 0.04fF
C1573 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C1574 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# gnd 0.05fF
C1575 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/a_n5_n50# gnd 0.05fF
C1576 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# 0.08fF
C1577 multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# 0.04fF
C1578 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.46fF
C1579 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C1580 gnd multiplier_0/and_7/nand_0/a_n5_n50# 0.05fF
C1581 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/m1_n2858_385# 0.20fF
C1582 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.13fF
C1583 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_1/m1_n1726_385# 0.20fF
C1584 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# gnd 0.11fF
C1585 multiplier_0/4bitadder_1/fulladder_0/m1_411_129# vdd 0.79fF
C1586 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1587 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# 0.13fF
C1588 gnd multiplier_0/and_0/nand_0/a_n5_n50# 0.05fF
C1589 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C1590 multiplier_0/and_9/inverter_0/w_0_0# multiplier_0/and_9/m1_59_58# 0.08fF
C1591 inA2 multiplier_0/and_6/m1_59_58# 0.20fF
C1592 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# 0.13fF
C1593 inA2 multiplier_0/and_10/m1_59_58# 0.20fF
C1594 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# 0.13fF
C1595 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C1596 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# 0.63fF
C1597 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# vdd 0.13fF
C1598 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# multiplier_0/m1_n611_n78# 0.08fF
C1599 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# gnd 0.13fF
C1600 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# vdd 0.04fF
C1601 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# 0.08fF
C1602 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/m1_411_129# 0.13fF
C1603 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C1604 multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/a_n5_n50# gnd 0.05fF
C1605 vdd multiplier_0/m1_n2157_n115# 2.94fF
C1606 inA1 inA2 1.92fF
C1607 multiplier_0/and_1/m1_59_58# multiplier_0/m1_n294_n107# 0.03fF
C1608 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/w_n27_n3# multiplier_0/m1_n294_n107# 0.13fF
C1609 multiplier_0/and_13/nand_0/w_n27_n3# inB3 0.13fF
C1610 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n3602_n1349# 0.13fF
C1611 multiplier_0/m1_n2288_n756# multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# 0.20fF
C1612 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# 0.08fF
C1613 multiplier_0/4bitadder_0/fulladder_1/m1_411_129# vdd 0.79fF
C1614 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# gnd 0.13fF
C1615 multiplier_0/m1_n4235_n2059# multiplier_0/m1_n4992_n2575# 3.96fF
C1616 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# gnd 0.23fF
C1617 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# 0.13fF
C1618 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# P5 0.20fF
C1619 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# vdd 0.10fF
C1620 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# 0.03fF
C1621 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/a_n5_n50# 0.08fF
C1622 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/w_n27_n3# multiplier_0/m1_n1820_n104# 0.13fF
C1623 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# 0.03fF
C1624 inA2 inB3 1.16fF
C1625 gnd multiplier_0/and_6/m1_59_58# 0.07fF
C1626 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# 0.08fF
C1627 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/w_n27_n3# vdd 0.04fF
C1628 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# vdd 0.10fF
C1629 multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# vdd 0.10fF
C1630 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# 0.13fF
C1631 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# gnd 0.05fF
C1632 multiplier_0/and_10/inverter_0/w_0_0# multiplier_0/m1_n3306_n1348# 0.04fF
C1633 gnd multiplier_0/and_10/m1_59_58# 0.07fF
C1634 multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_1/w_0_0# vdd 0.13fF
C1635 multiplier_0/m1_n2688_n2050# multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# 0.08fF
C1636 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# 0.08fF
C1637 gnd inA1 0.33fF
C1638 multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_0/w_0_0# 0.08fF
C1639 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# multiplier_0/m1_n4992_n2575# 0.13fF
C1640 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# gnd 0.11fF
C1641 multiplier_0/m1_n1128_n767# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# 0.20fF
C1642 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C1643 gnd multiplier_0/and_15/m1_59_58# 0.07fF
C1644 vdd multiplier_0/and_5/nand_0/w_n27_n3# 0.04fF
C1645 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# vdd 0.10fF
C1646 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# 0.30fF
C1647 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# multiplier_0/m1_n4992_n2575# 0.32fF
C1648 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# 0.13fF
C1649 multiplier_0/m1_n3416_n801# multiplier_0/m1_n3306_n1348# 0.26fF
C1650 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# gnd 0.23fF
C1651 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# 0.13fF
C1652 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# vdd 0.04fF
C1653 inB1 multiplier_0/and_6/nand_0/w_n27_n3# 0.13fF
C1654 multiplier_0/m1_n4235_n2059# vdd 1.21fF
C1655 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# vdd 0.04fF
C1656 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/w_n27_n3# multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# 0.13fF
C1657 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# multiplier_0/4bitadder_2/m1_n594_383# 0.13fF
C1658 multiplier_0/m1_n3849_n2792# Gnd 14.99fF
C1659 multiplier_0/and_15/m1_59_58# Gnd 0.67fF
C1660 multiplier_0/and_15/inverter_0/w_0_0# Gnd 0.73fF
C1661 multiplier_0/and_15/nand_0/a_n5_n50# Gnd 0.02fF
C1662 inB3 Gnd 31.52fF
C1663 multiplier_0/and_15/nand_0/w_n27_n3# Gnd 1.55fF
C1664 multiplier_0/m1_n4201_n2800# Gnd 14.88fF
C1665 multiplier_0/and_14/m1_59_58# Gnd 0.67fF
C1666 multiplier_0/and_14/inverter_0/w_0_0# Gnd 0.73fF
C1667 multiplier_0/and_14/nand_0/a_n5_n50# Gnd 0.02fF
C1668 multiplier_0/and_14/nand_0/w_n27_n3# Gnd 1.55fF
C1669 multiplier_0/m1_n4533_n2563# Gnd 5.05fF
C1670 multiplier_0/and_13/m1_59_58# Gnd 0.67fF
C1671 multiplier_0/and_13/inverter_0/w_0_0# Gnd 0.73fF
C1672 multiplier_0/and_13/nand_0/a_n5_n50# Gnd 0.02fF
C1673 multiplier_0/and_13/nand_0/w_n27_n3# Gnd 1.55fF
C1674 multiplier_0/m1_n4992_n2575# Gnd 10.71fF
C1675 multiplier_0/and_12/m1_59_58# Gnd 0.67fF
C1676 multiplier_0/and_12/inverter_0/w_0_0# Gnd 0.73fF
C1677 multiplier_0/and_12/nand_0/a_n5_n50# Gnd 0.02fF
C1678 multiplier_0/and_12/nand_0/w_n27_n3# Gnd 1.55fF
C1679 multiplier_0/m1_n3602_n1349# Gnd 13.30fF
C1680 multiplier_0/and_11/m1_59_58# Gnd 0.67fF
C1681 multiplier_0/and_11/inverter_0/w_0_0# Gnd 0.73fF
C1682 multiplier_0/and_11/nand_0/a_n5_n50# Gnd 0.02fF
C1683 multiplier_0/and_11/nand_0/w_n27_n3# Gnd 1.55fF
C1684 multiplier_0/m1_n3306_n1348# Gnd 5.39fF
C1685 multiplier_0/and_10/m1_59_58# Gnd 0.67fF
C1686 multiplier_0/and_10/inverter_0/w_0_0# Gnd 0.73fF
C1687 multiplier_0/and_10/nand_0/a_n5_n50# Gnd 0.02fF
C1688 multiplier_0/and_10/nand_0/w_n27_n3# Gnd 1.55fF
C1689 multiplier_0/m1_n2968_n1347# Gnd 15.41fF
C1690 multiplier_0/and_9/m1_59_58# Gnd 0.67fF
C1691 multiplier_0/and_9/inverter_0/w_0_0# Gnd 0.73fF
C1692 multiplier_0/and_9/nand_0/a_n5_n50# Gnd 0.02fF
C1693 multiplier_0/and_9/nand_0/w_n27_n3# Gnd 1.55fF
C1694 multiplier_0/m1_n2617_n1342# Gnd 17.60fF
C1695 multiplier_0/and_8/m1_59_58# Gnd 0.67fF
C1696 multiplier_0/and_8/inverter_0/w_0_0# Gnd 0.73fF
C1697 multiplier_0/and_8/nand_0/a_n5_n50# Gnd 0.02fF
C1698 inB2 Gnd 42.48fF
C1699 multiplier_0/and_8/nand_0/w_n27_n3# Gnd 1.55fF
C1700 multiplier_0/m1_n2782_n115# Gnd 13.78fF
C1701 multiplier_0/and_7/m1_59_58# Gnd 0.67fF
C1702 multiplier_0/and_7/inverter_0/w_0_0# Gnd 0.73fF
C1703 multiplier_0/and_7/nand_0/a_n5_n50# Gnd 0.02fF
C1704 multiplier_0/and_7/nand_0/w_n27_n3# Gnd 1.55fF
C1705 multiplier_0/m1_n2469_n98# Gnd 5.23fF
C1706 multiplier_0/and_6/m1_59_58# Gnd 0.67fF
C1707 multiplier_0/and_6/inverter_0/w_0_0# Gnd 0.73fF
C1708 multiplier_0/and_6/nand_0/a_n5_n50# Gnd 0.02fF
C1709 multiplier_0/and_6/nand_0/w_n27_n3# Gnd 1.55fF
C1710 multiplier_0/m1_n2157_n115# Gnd 15.60fF
C1711 multiplier_0/and_5/m1_59_58# Gnd 0.67fF
C1712 multiplier_0/and_5/inverter_0/w_0_0# Gnd 0.73fF
C1713 multiplier_0/and_5/nand_0/a_n5_n50# Gnd 0.02fF
C1714 multiplier_0/and_5/nand_0/w_n27_n3# Gnd 1.55fF
C1715 multiplier_0/m1_n1820_n104# Gnd 17.35fF
C1716 multiplier_0/and_4/m1_59_58# Gnd 0.67fF
C1717 multiplier_0/and_4/inverter_0/w_0_0# Gnd 0.73fF
C1718 multiplier_0/and_4/nand_0/a_n5_n50# Gnd 0.02fF
C1719 inB1 Gnd 3.05fF
C1720 multiplier_0/and_4/nand_0/w_n27_n3# Gnd 1.55fF
C1721 multiplier_0/m1_n980_n67# Gnd 12.07fF
C1722 multiplier_0/and_3/m1_59_58# Gnd 0.67fF
C1723 multiplier_0/and_3/inverter_0/w_0_0# Gnd 0.73fF
C1724 multiplier_0/and_3/nand_0/a_n5_n50# Gnd 0.02fF
C1725 inA3 Gnd 160.12fF
C1726 multiplier_0/and_3/nand_0/w_n27_n3# Gnd 1.55fF
C1727 multiplier_0/m1_n611_n78# Gnd 4.18fF
C1728 multiplier_0/and_2/m1_59_58# Gnd 0.67fF
C1729 multiplier_0/and_2/inverter_0/w_0_0# Gnd 0.73fF
C1730 multiplier_0/and_2/nand_0/a_n5_n50# Gnd 0.02fF
C1731 inA2 Gnd 158.53fF
C1732 multiplier_0/and_2/nand_0/w_n27_n3# Gnd 1.55fF
C1733 multiplier_0/m1_n294_n107# Gnd 2.52fF
C1734 multiplier_0/and_1/m1_59_58# Gnd 0.67fF
C1735 multiplier_0/and_1/inverter_0/w_0_0# Gnd 0.73fF
C1736 multiplier_0/and_1/nand_0/a_n5_n50# Gnd 0.02fF
C1737 inA1 Gnd 152.35fF
C1738 multiplier_0/and_1/nand_0/w_n27_n3# Gnd 1.55fF
C1739 gnd Gnd 892.94fF
C1740 P0 Gnd 63.22fF
C1741 vdd Gnd 854.43fF
C1742 multiplier_0/and_0/m1_59_58# Gnd 0.67fF
C1743 multiplier_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1744 multiplier_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1745 inA0 Gnd 150.49fF
C1746 inB0 Gnd 39.24fF
C1747 multiplier_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1748 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1749 P3 Gnd 11.64fF
C1750 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C1751 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C1752 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1753 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1754 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1755 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1756 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1757 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1758 multiplier_0/4bitadder_2/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C1759 multiplier_0/4bitadder_2/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1760 multiplier_0/4bitadder_2/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C1761 multiplier_0/4bitadder_2/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1762 multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1763 multiplier_0/4bitadder_2/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1764 multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_1/w_0_0# Gnd 0.73fF
C1765 multiplier_0/4bitadder_2/fulladder_2/m1_n28_112# Gnd 0.55fF
C1766 multiplier_0/4bitadder_2/fulladder_2/or_0/inverter_0/w_0_0# Gnd 0.73fF
C1767 multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/a_n5_n50# Gnd 0.02fF
C1768 P7 Gnd 18.05fF
C1769 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n44# Gnd 0.68fF
C1770 multiplier_0/4bitadder_2/fulladder_2/or_0/m1_38_n14# Gnd 0.69fF
C1771 multiplier_0/4bitadder_2/fulladder_2/or_0/nand_0/w_n27_n3# Gnd 1.55fF
C1772 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1773 P6 Gnd 7.67fF
C1774 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_140_2# Gnd 1.13fF
C1775 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_144_120# Gnd 1.16fF
C1776 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1777 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1778 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1779 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1780 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1781 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1782 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/m1_51_58# Gnd 1.80fF
C1783 multiplier_0/4bitadder_2/fulladder_2/m1_411_129# Gnd 3.30fF
C1784 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1785 multiplier_0/4bitadder_2/fulladder_2/m1_n30_n19# Gnd 4.57fF
C1786 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/m1_59_58# Gnd 0.67fF
C1787 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1788 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1789 multiplier_0/4bitadder_2/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1790 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1791 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C1792 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C1793 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1794 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1795 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1796 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1797 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1798 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1799 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C1800 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1801 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C1802 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1803 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1804 multiplier_0/4bitadder_2/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1805 multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_1/w_0_0# Gnd 0.73fF
C1806 multiplier_0/4bitadder_2/fulladder_1/m1_n28_112# Gnd 0.55fF
C1807 multiplier_0/4bitadder_2/fulladder_1/or_0/inverter_0/w_0_0# Gnd 0.73fF
C1808 multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/a_n5_n50# Gnd 0.02fF
C1809 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n44# Gnd 0.68fF
C1810 multiplier_0/4bitadder_2/fulladder_1/or_0/m1_38_n14# Gnd 0.69fF
C1811 multiplier_0/4bitadder_2/fulladder_1/or_0/nand_0/w_n27_n3# Gnd 1.55fF
C1812 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1813 P5 Gnd 10.79fF
C1814 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_140_2# Gnd 1.13fF
C1815 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_144_120# Gnd 1.16fF
C1816 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1817 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1818 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1819 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1820 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1821 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1822 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/m1_51_58# Gnd 1.80fF
C1823 multiplier_0/4bitadder_2/fulladder_1/m1_411_129# Gnd 3.30fF
C1824 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1825 multiplier_0/4bitadder_2/fulladder_1/m1_n30_n19# Gnd 4.57fF
C1826 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/m1_59_58# Gnd 0.67fF
C1827 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1828 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1829 multiplier_0/4bitadder_2/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1830 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1831 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C1832 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C1833 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1834 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1835 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1836 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1837 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1838 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1839 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C1840 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1841 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C1842 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1843 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1844 multiplier_0/4bitadder_2/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1845 multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_1/w_0_0# Gnd 0.73fF
C1846 multiplier_0/4bitadder_2/fulladder_0/m1_n28_112# Gnd 0.55fF
C1847 multiplier_0/4bitadder_2/fulladder_0/or_0/inverter_0/w_0_0# Gnd 0.73fF
C1848 multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/a_n5_n50# Gnd 0.02fF
C1849 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n44# Gnd 0.68fF
C1850 multiplier_0/4bitadder_2/fulladder_0/or_0/m1_38_n14# Gnd 0.69fF
C1851 multiplier_0/4bitadder_2/fulladder_0/or_0/nand_0/w_n27_n3# Gnd 1.55fF
C1852 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1853 P4 Gnd 17.15fF
C1854 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_140_2# Gnd 1.13fF
C1855 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_144_120# Gnd 1.16fF
C1856 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1857 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1858 multiplier_0/4bitadder_2/m1_n594_383# Gnd 3.77fF
C1859 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1860 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1861 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1862 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1863 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/m1_51_58# Gnd 1.80fF
C1864 multiplier_0/4bitadder_2/fulladder_0/m1_411_129# Gnd 3.30fF
C1865 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1866 multiplier_0/4bitadder_2/fulladder_0/m1_n30_n19# Gnd 4.57fF
C1867 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/m1_59_58# Gnd 0.67fF
C1868 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1869 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1870 multiplier_0/4bitadder_2/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1871 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1872 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C1873 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C1874 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1875 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1876 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1877 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1878 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1879 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1880 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C1881 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1882 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C1883 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1884 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1885 multiplier_0/4bitadder_2/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1886 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1887 P2 Gnd 33.73fF
C1888 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C1889 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C1890 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1891 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1892 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1893 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1894 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1895 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1896 multiplier_0/4bitadder_1/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C1897 multiplier_0/4bitadder_1/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1898 multiplier_0/4bitadder_1/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C1899 multiplier_0/4bitadder_1/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1900 multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1901 multiplier_0/4bitadder_1/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1902 multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_1/w_0_0# Gnd 0.73fF
C1903 multiplier_0/4bitadder_1/fulladder_2/m1_n28_112# Gnd 0.55fF
C1904 multiplier_0/4bitadder_1/fulladder_2/or_0/inverter_0/w_0_0# Gnd 0.73fF
C1905 multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/a_n5_n50# Gnd 0.02fF
C1906 multiplier_0/m1_n4235_n2059# Gnd 23.75fF
C1907 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n44# Gnd 0.68fF
C1908 multiplier_0/4bitadder_1/fulladder_2/or_0/m1_38_n14# Gnd 0.69fF
C1909 multiplier_0/4bitadder_1/fulladder_2/or_0/nand_0/w_n27_n3# Gnd 1.55fF
C1910 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1911 multiplier_0/m1_n3123_n2056# Gnd 14.01fF
C1912 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_140_2# Gnd 1.13fF
C1913 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_144_120# Gnd 1.16fF
C1914 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1915 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1916 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1917 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1918 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1919 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1920 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/m1_51_58# Gnd 1.80fF
C1921 multiplier_0/4bitadder_1/fulladder_2/m1_411_129# Gnd 3.30fF
C1922 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1923 multiplier_0/4bitadder_1/fulladder_2/m1_n30_n19# Gnd 4.57fF
C1924 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/m1_59_58# Gnd 0.67fF
C1925 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1926 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1927 multiplier_0/4bitadder_1/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1928 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1929 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C1930 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C1931 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1932 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1933 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1934 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1935 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1936 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1937 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C1938 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1939 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C1940 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1941 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1942 multiplier_0/4bitadder_1/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1943 multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_1/w_0_0# Gnd 0.73fF
C1944 multiplier_0/4bitadder_1/fulladder_1/m1_n28_112# Gnd 0.55fF
C1945 multiplier_0/4bitadder_1/fulladder_1/or_0/inverter_0/w_0_0# Gnd 0.73fF
C1946 multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/a_n5_n50# Gnd 0.02fF
C1947 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n44# Gnd 0.68fF
C1948 multiplier_0/4bitadder_1/fulladder_1/or_0/m1_38_n14# Gnd 0.69fF
C1949 multiplier_0/4bitadder_1/fulladder_1/or_0/nand_0/w_n27_n3# Gnd 1.55fF
C1950 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1951 multiplier_0/m1_n2688_n2050# Gnd 12.97fF
C1952 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_140_2# Gnd 1.13fF
C1953 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_144_120# Gnd 1.16fF
C1954 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1955 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1956 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1957 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1958 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1959 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1960 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/m1_51_58# Gnd 1.80fF
C1961 multiplier_0/4bitadder_1/fulladder_1/m1_411_129# Gnd 3.30fF
C1962 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1963 multiplier_0/4bitadder_1/fulladder_1/m1_n30_n19# Gnd 4.57fF
C1964 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/m1_59_58# Gnd 0.67fF
C1965 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1966 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1967 multiplier_0/4bitadder_1/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1968 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1969 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C1970 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C1971 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1972 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1973 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1974 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1975 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C1976 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C1977 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C1978 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C1979 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C1980 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C1981 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C1982 multiplier_0/4bitadder_1/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C1983 multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_1/w_0_0# Gnd 0.73fF
C1984 multiplier_0/4bitadder_1/fulladder_0/m1_n28_112# Gnd 0.55fF
C1985 multiplier_0/4bitadder_1/fulladder_0/or_0/inverter_0/w_0_0# Gnd 0.73fF
C1986 multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/a_n5_n50# Gnd 0.02fF
C1987 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n44# Gnd 0.68fF
C1988 multiplier_0/4bitadder_1/fulladder_0/or_0/m1_38_n14# Gnd 0.69fF
C1989 multiplier_0/4bitadder_1/fulladder_0/or_0/nand_0/w_n27_n3# Gnd 1.55fF
C1990 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C1991 multiplier_0/m1_n2369_n2126# Gnd 29.97fF
C1992 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_140_2# Gnd 1.13fF
C1993 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_144_120# Gnd 1.16fF
C1994 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C1995 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C1996 multiplier_0/4bitadder_1/m1_n594_383# Gnd 3.77fF
C1997 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C1998 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C1999 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C2000 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C2001 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/m1_51_58# Gnd 1.80fF
C2002 multiplier_0/4bitadder_1/fulladder_0/m1_411_129# Gnd 3.30fF
C2003 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C2004 multiplier_0/4bitadder_1/fulladder_0/m1_n30_n19# Gnd 4.57fF
C2005 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/m1_59_58# Gnd 0.67fF
C2006 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# Gnd 0.73fF
C2007 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C2008 multiplier_0/4bitadder_1/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C2009 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C2010 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C2011 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C2012 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C2013 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C2014 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C2015 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C2016 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C2017 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C2018 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C2019 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C2020 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C2021 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C2022 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C2023 multiplier_0/4bitadder_1/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C2024 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C2025 P1 Gnd 51.61fF
C2026 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C2027 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C2028 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C2029 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C2030 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C2031 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C2032 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C2033 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C2034 multiplier_0/4bitadder_0/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C2035 multiplier_0/4bitadder_0/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C2036 multiplier_0/4bitadder_0/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C2037 multiplier_0/4bitadder_0/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C2038 multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C2039 multiplier_0/4bitadder_0/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C2040 multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_1/w_0_0# Gnd 0.73fF
C2041 multiplier_0/4bitadder_0/fulladder_2/m1_n28_112# Gnd 0.55fF
C2042 multiplier_0/4bitadder_0/fulladder_2/or_0/inverter_0/w_0_0# Gnd 0.73fF
C2043 multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/a_n5_n50# Gnd 0.02fF
C2044 multiplier_0/m1_n3416_n801# Gnd 24.93fF
C2045 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n44# Gnd 0.68fF
C2046 multiplier_0/4bitadder_0/fulladder_2/or_0/m1_38_n14# Gnd 0.69fF
C2047 multiplier_0/4bitadder_0/fulladder_2/or_0/nand_0/w_n27_n3# Gnd 1.55fF
C2048 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C2049 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_140_2# Gnd 1.13fF
C2050 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_144_120# Gnd 1.16fF
C2051 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C2052 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C2053 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C2054 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C2055 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C2056 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C2057 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/m1_51_58# Gnd 1.80fF
C2058 multiplier_0/4bitadder_0/fulladder_2/m1_411_129# Gnd 3.30fF
C2059 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C2060 multiplier_0/4bitadder_0/fulladder_2/m1_n30_n19# Gnd 4.57fF
C2061 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/m1_59_58# Gnd 0.67fF
C2062 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/inverter_0/w_0_0# Gnd 0.73fF
C2063 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C2064 multiplier_0/4bitadder_0/fulladder_2/halfadder_1/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C2065 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C2066 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C2067 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C2068 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C2069 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C2070 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C2071 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C2072 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C2073 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C2074 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C2075 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C2076 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C2077 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C2078 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C2079 multiplier_0/4bitadder_0/fulladder_2/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C2080 multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_1/w_0_0# Gnd 0.73fF
C2081 multiplier_0/4bitadder_0/fulladder_1/m1_n28_112# Gnd 0.55fF
C2082 multiplier_0/4bitadder_0/fulladder_1/or_0/inverter_0/w_0_0# Gnd 0.73fF
C2083 multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/a_n5_n50# Gnd 0.02fF
C2084 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n44# Gnd 0.68fF
C2085 multiplier_0/4bitadder_0/fulladder_1/or_0/m1_38_n14# Gnd 0.69fF
C2086 multiplier_0/4bitadder_0/fulladder_1/or_0/nand_0/w_n27_n3# Gnd 1.55fF
C2087 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C2088 multiplier_0/m1_n1473_n1361# Gnd 2.52fF
C2089 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_140_2# Gnd 1.13fF
C2090 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_144_120# Gnd 1.16fF
C2091 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C2092 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C2093 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C2094 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C2095 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C2096 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C2097 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/m1_51_58# Gnd 1.80fF
C2098 multiplier_0/4bitadder_0/fulladder_1/m1_411_129# Gnd 3.30fF
C2099 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C2100 multiplier_0/4bitadder_0/fulladder_1/m1_n30_n19# Gnd 4.57fF
C2101 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/m1_59_58# Gnd 0.67fF
C2102 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/inverter_0/w_0_0# Gnd 0.73fF
C2103 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C2104 multiplier_0/4bitadder_0/fulladder_1/halfadder_1/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C2105 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C2106 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C2107 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C2108 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C2109 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C2110 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C2111 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C2112 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C2113 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C2114 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C2115 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C2116 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C2117 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C2118 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C2119 multiplier_0/4bitadder_0/fulladder_1/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C2120 multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_1/w_0_0# Gnd 0.73fF
C2121 multiplier_0/4bitadder_0/fulladder_0/m1_n28_112# Gnd 0.55fF
C2122 multiplier_0/4bitadder_0/fulladder_0/or_0/inverter_0/w_0_0# Gnd 0.73fF
C2123 multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/a_n5_n50# Gnd 0.02fF
C2124 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n44# Gnd 0.68fF
C2125 multiplier_0/4bitadder_0/fulladder_0/or_0/m1_38_n14# Gnd 0.69fF
C2126 multiplier_0/4bitadder_0/fulladder_0/or_0/nand_0/w_n27_n3# Gnd 1.55fF
C2127 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C2128 multiplier_0/m1_n1128_n767# Gnd 24.10fF
C2129 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_140_2# Gnd 1.13fF
C2130 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_144_120# Gnd 1.16fF
C2131 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C2132 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C2133 multiplier_0/4bitadder_0/m1_n594_383# Gnd 3.77fF
C2134 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C2135 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C2136 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C2137 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C2138 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/m1_51_58# Gnd 1.80fF
C2139 multiplier_0/4bitadder_0/fulladder_0/m1_411_129# Gnd 3.30fF
C2140 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C2141 multiplier_0/4bitadder_0/fulladder_0/m1_n30_n19# Gnd 4.57fF
C2142 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/m1_59_58# Gnd 0.67fF
C2143 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/inverter_0/w_0_0# Gnd 0.73fF
C2144 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C2145 multiplier_0/4bitadder_0/fulladder_0/halfadder_1/and_0/nand_0/w_n27_n3# Gnd 1.55fF
C2146 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/a_n5_n50# Gnd 0.02fF
C2147 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_140_2# Gnd 1.13fF
C2148 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_144_120# Gnd 1.16fF
C2149 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_3/w_n27_n3# Gnd 1.55fF
C2150 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/a_n5_n50# Gnd 0.02fF
C2151 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_2/w_n27_n3# Gnd 1.55fF
C2152 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/a_n5_n50# Gnd 0.02fF
C2153 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_0/w_n27_n3# Gnd 1.55fF
C2154 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/a_n5_n50# Gnd 0.02fF
C2155 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/m1_51_58# Gnd 1.80fF
C2156 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/xor_0/nand_1/w_n27_n3# Gnd 1.55fF
C2157 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/m1_59_58# Gnd 0.67fF
C2158 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/inverter_0/w_0_0# Gnd 0.73fF
C2159 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/a_n5_n50# Gnd 0.02fF
C2160 multiplier_0/4bitadder_0/fulladder_0/halfadder_0/and_0/nand_0/w_n27_n3# Gnd 1.55fF

Vd0 P7 gnd DC 0V


.tran 0.1n 40n

* for P0
.measure tran td_0_lh TRIG v(inA2) VAL=0.5 FALL=2 TARG v(P0) val=0.5 RISE=2
.measure tran td_0_hl TRIG v(inA2) VAL=0.5 RISE=2 TARG v(P0) val=0.5 FALL=2

* for P1
.measure tran td_1_lh TRIG v(inA2) VAL=0.5 FALL=2 TARG v(P1) val=0.5 RISE=2
.measure tran td_1_hl TRIG v(inA2) VAL=0.5 RISE=2 TARG v(P1) val=0.5 FALL=2

* for P2
.measure tran td_2_lh TRIG v(inA2) VAL=0.5 RISE=1 TARG v(P2) val=0.5 RISE=1
.measure tran td_2_hl TRIG v(inA2) VAL=0.5 FALL=2 TARG v(P2) val=0.5 FALL=2


* for P3
.measure tran td_3_lh TRIG v(inA2) VAL=0.5 RISE=1 TARG v(P3) val=0.5 RISE=1
.measure tran td_3_hl TRIG v(inA2) VAL=0.5 FALL=2 TARG v(P3) val=0.5 FALL=2


* for P4
.measure tran td_4_lh TRIG v(inA2) VAL=0.5 RISE=1 TARG v(P4) val=0.5 RISE=1
.measure tran td_4_hl TRIG v(inA2) VAL=0.5 FALL=2 TARG v(P4) val=0.5 FALL=2


* for P5
.measure tran td_5_lh TRIG v(inA2) VAL=0.5 FALL=2 TARG v(P5) val=0.5 RISE=2
.measure tran td_5_hl TRIG v(inA2) VAL=0.5 RISE=2 TARG v(P5) val=0.5 FALL=2

* for P6
.measure tran td_6_lh TRIG v(inA2) VAL=0.5 FALL=2 TARG v(P6) val=0.5 RISE=2
.measure tran td_6_hl TRIG v(inA2) VAL=0.5 RISE=2 TARG v(P6) val=0.5 FALL=2

* for P7
.measure tran td_7_lh TRIG v(inA2) VAL=0.5 RISE=1 TARG v(P7) val=0.5 RISE=1
.measure tran td_7_hl TRIG v(inA2) VAL=0.5 FALL=2 TARG v(P7) val=0.5 FALL=2


.control
* set hcopycolor = 1
* set color0=white
* set color1=black

run
plot v(inA0) v(inA1)+10 v(inA2)+20 v(inA3)+30
plot v(inB0) v(inB1)+10 v(inB2)+20 v(inB3)+30

plot v(P0) v(P1)+10 v(P2)+20 v(P3)+30 v(P4)+40 v(P5)+50 v(P6)+60 v(P7)+70

plot Vd0#branch

.endc

* .measure tran idt INTEG i(Vd0) from=0 to=20n

.end