magic
tech scmos
timestamp 1669292255
<< metal1 >>
rect -4 95 3 99
rect 122 69 126 77
rect -4 29 3 33
<< metal2 >>
rect 53 136 60 140
rect 57 -2 64 2
use or  or_0
timestamp 1669292154
transform 1 0 9 0 1 75
box -9 -75 115 63
<< labels >>
rlabel metal1 -4 29 3 33 3 inB
rlabel metal1 -4 95 3 99 3 inA
rlabel metal2 53 136 60 140 5 vdd
rlabel metal2 57 -2 64 2 1 gnd
rlabel metal1 122 69 126 77 7 out
<< end >>
