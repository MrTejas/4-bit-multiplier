magic
tech scmos
timestamp 1669286840
<< nwell >>
rect -27 -3 30 24
<< ntransistor >>
rect -9 -50 -5 -42
rect 6 -50 10 -42
<< ptransistor >>
rect -9 8 -5 17
rect 6 8 10 17
<< ndiffusion >>
rect -13 -50 -9 -42
rect -5 -50 -4 -42
rect 4 -50 6 -42
rect 10 -50 13 -42
<< pdiffusion >>
rect -12 8 -9 17
rect -5 8 -4 17
rect 4 8 6 17
rect 10 8 13 17
<< ndcontact >>
rect -21 -50 -13 -42
rect -4 -50 4 -42
rect 13 -50 21 -42
<< pdcontact >>
rect -20 8 -12 17
rect -4 8 4 17
rect 13 8 21 17
<< polysilicon >>
rect -9 17 -5 20
rect 6 17 10 20
rect -9 -25 -5 8
rect -9 -42 -5 -29
rect 6 -34 10 8
rect 6 -42 10 -38
rect -9 -54 -5 -50
rect 6 -54 10 -50
<< polycontact >>
rect -9 -29 -5 -25
rect 6 -38 10 -34
<< metal1 >>
rect -27 26 30 32
rect -4 17 4 26
rect -20 -14 -12 8
rect 13 -13 21 8
rect 13 -14 30 -13
rect -20 -21 30 -14
rect -28 -29 -9 -25
rect -28 -38 6 -34
rect 13 -42 21 -21
rect -21 -57 -13 -50
rect -28 -64 26 -57
<< end >>
