* SPICE3 file created from nand_test.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY=5
.option scale=0.09u
.global vdd gnd


Vdd vdd gnd 'SUPPLY'
vinA inA gnd pulse 0 'SUPPLY' 0ns 0.1ns 0.1ns 10ns 20ns
vinB inB gnd pulse 0 'SUPPLY' 0ns 0.1ns 0.1ns 20ns 40ns



M1000 out inB nand_0/a_n5_n50# Gnd nfet w=8 l=4
+  ad=88 pd=38 as=88 ps=38
M1001 nand_0/a_n5_n50# inA gnd Gnd nfet w=8 l=4
+  ad=0 pd=0 as=96 ps=40
M1002 out inB vdd nand_0/w_n27_n3# pfet w=9 l=4
+  ad=198 pd=80 as=99 ps=40
M1003 vdd inA out nand_0/w_n27_n3# pfet w=9 l=4
+  ad=0 pd=0 as=0 ps=0
C0 out inA 0.24fF
C1 inB gnd 0.11fF
C2 inB out 0.20fF
C3 inB nand_0/a_n5_n50# 0.11fF
C4 vdd nand_0/w_n27_n3# 0.04fF
C5 nand_0/w_n27_n3# inA 0.13fF
C6 inB nand_0/w_n27_n3# 0.13fF
C7 inB inA 0.48fF
C8 out nand_0/w_n27_n3# 0.13fF


.tran 0.1n 40n

.control
* set hcopycolor = 1
* set color0=white
* set color1=black

run
plot v(inA) 10+v(inB) v(out)+20

.endc

.end