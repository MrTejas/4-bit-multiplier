
.include 22nm_MGK.pm
.include and2.sub
.include halfadder.sub
.include fulladder.sub
.include 4bitadder.sub
.include multiplier.sub

.param SUPPLY = 1
.param LAMBDA = 22n 

*given lambda = length and length is given as 22nm thus lambda = 22nm

.param width_N =  {2*LAMBDA}
.param width_P =   {2*LAMBDA} 
.global gnd vdd

VDS vdd gnd DC 'SUPPLY'
* va A0 gnd pulse 0 1 0ns 10ps 10ps 10ns 20ns
* vb A1 gnd pulse 0 1 10ns 10ps 10ps 10ns 20ns
* vc A2 gnd pulse 0 1 0ns 10ps 10ps 10ns 20ns
* vd A3 gnd pulse 0 1 10ns 10ps 10ps 10ns 20ns

* ve B0 gnd pulse 0 1 0ns 10ps 10ps 10ns 20ns
* vf B1 gnd pulse 0 1 0ns 10ps 10ps 10ns 20ns
* vg B2 gnd pulse 0 1 0ns 10ps 10ps 10ns 20ns
* vh B3 gnd pulse 0 1 0ns 10ps 10ps 10ns 20ns

* va A0 gnd 1 DC
* vl A1 gnd 1 DC
* vp A2 gnd 1 DC
* vk A3 gnd 1 DC

* vj B0 gnd 1 DC
* vd B1 gnd 1 DC
* vg B2 gnd 1 DC
* vf B3 gnd 1 DC

va A0 gnd 0 DC
vb A1 gnd 'SUPPLY' DC
vc A2 gnd pulse 1 0 0ns 10ps 10ps 10ns 20ns
vd A3 gnd 0 DC

ve B0 gnd pulse 0 1 0ns 10ps 10ps 10ns 20ns
vf B1 gnd pulse 0 1 0ns 10ps 10ps 10ns 20ns
vg B2 gnd pulse 1 0 0ns 10ps 10ps 10ns 20ns
vh B3 gnd 0 DC

* X1 A0 B0 S0 C1 gnd high HalfAdder
* X2 A1 B1 C1 S1 C2 gnd high FullAdder
* X3 A2 B2 C2 S2 C3 gnd high FullAdder
* X4 A3 B3 C3 S3 C4 gnd high FullAdder

X1 A0 A1 A2 A3 B0 B1 B2 B3 P0 P1 P2 P3 P4 P5 P6 P7 gnd vdd multiplier

Vd0 P7 gnd DC 0V

.tran 1n 120n

* for P0
.measure tran td_0_lh TRIG v(A2) VAL=0.5 FALL=2 TARG v(P0) val=0.5 RISE=2
.measure tran td_0_hl TRIG v(A2) VAL=0.5 RISE=2 TARG v(P0) val=0.5 FALL=2

* for P1
.measure tran td_1_lh TRIG v(A2) VAL=0.5 FALL=2 TARG v(P1) val=0.5 RISE=2
.measure tran td_1_hl TRIG v(A2) VAL=0.5 RISE=2 TARG v(P1) val=0.5 FALL=2

* for P2
.measure tran td_2_lh TRIG v(A2) VAL=0.5 FALL=2 TARG v(P2) val=0.5 RISE=2
.measure tran td_2_hl TRIG v(A2) VAL=0.5 RISE=2 TARG v(P2) val=0.5 FALL=2


* for P3
.measure tran td_3_lh TRIG v(A2) VAL=0.5 RISE=1 TARG v(P3) val=0.5 RISE=1
.measure tran td_3_hl TRIG v(A2) VAL=0.5 FALL=2 TARG v(P3) val=0.5 FALL=2


* for P4
.measure tran td_4_lh TRIG v(A2) VAL=0.5 RISE=1 TARG v(P4) val=0.5 RISE=1
.measure tran td_4_hl TRIG v(A2) VAL=0.5 FALL=2 TARG v(P4) val=0.5 FALL=2


* for P5
.measure tran td_5_lh TRIG v(A2) VAL=0.5 FALL=2 TARG v(P5) val=0.5 RISE=2
.measure tran td_5_hl TRIG v(A2) VAL=0.5 RISE=2 TARG v(P5) val=0.5 FALL=2

* for P6
.measure tran td_6_lh TRIG v(A2) VAL=0.5 FALL=2 TARG v(P6) val=0.5 RISE=2
.measure tran td_6_hl TRIG v(A2) VAL=0.5 RISE=2 TARG v(P6) val=0.5 FALL=2

* for P7
.measure tran td_7_lh TRIG v(A2) VAL=0.5 RISE=1 TARG v(P7) val=0.5 RISE=1
.measure tran td_7_hl TRIG v(A2) VAL=0.5 FALL=2 TARG v(P7) val=0.5 FALL=2


1

* .measure tran td7 TRIG v(A0) VAL=0.5 RISE=1 TARG v(P3) val=0.5 FALL=1
* .measure tran td3 TRIG v(A0) VAL=0.5 RISE=1 TARG v(P7) val=0.5 FALL=1

.control
run

tran 1n 120n
plot v(A0) 2+v(A1) 4+v(A2) 6+v(A3) 
plot v(B0) 2+v(B1) 4+v(B2) 6+v(B3) 
plot v(P0) 2+v(P1) 4+v(P2) 6+v(P3) 8+v(P4) 10+v(P5) 12+v(P6) 14+v(P7) 

plot Vd0#branch
.endc

* .measure tran idt INTEG i(Vd0) from=0 to=20n


.end