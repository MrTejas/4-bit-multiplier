4 bit multiplier Circuit
.include 22nm_MGK.pm
.param SUPPLY = 2
.global vdd gnd


* -----------------SUBCIRCUIT OF 2 input AND--------------
.subckt and2 a b y gnd

* .param SUPPLY = 0.6
.global vdd gnd
.param width_nmos=44
.param width_pmos=44
.param length_nmos=22
.param length_pmos=22

Vss1 vdd gnd DC 'SUPPLY'


Mp1 n1 a vdd vdd pmos W=44nm L=22nm
Mp2 n1 b vdd vdd pmos W=44nm L=22nm
Mp3 y n1 vdd vdd pmos W=44nm L=22nm

Mn1 n1 a n2 n2 nmos W=44nm L=22nm
Mn2 n2 b gnd gnd nmos W=44nm L=22nm
Mn3 y n1 gnd gnd nmos W=44nm L=22nm

.ends and2
* ----------------------END OF SUBCIRCUIT----------------------
.end


* -----------------SUBCIRCUIT OF 3-BIT FULL ADDER--------------
.subckt FullAdder a b c n_sum n_carry gnd

* .param SUPPLY = 0.6
.global vdd gnd
* .param width_nmos=44
* .param width_pmos=44
* .param length_nmos=22
* .param length_pmos=22

Vss2 vdd gnd DC 'SUPPLY'


Mp1     n0 a vdd vdd pmos W=44nm L=22nm
Mp2     n2 b n0  n0  pmos W=44nm L=22nm
Mp3     n3 a vdd vdd pmos W=44nm L=22nm
Mp4     n3 b vdd vdd pmos W=44nm L=22nm
Mp5     n2 c n3  n3  pmos W=44nm L=22nm
Mp6     n5 c vdd vdd pmos W=44nm L=22nm
Mp7     n5 a vdd vdd pmos W=44nm L=22nm
Mp8     n5 b vdd vdd pmos W=44nm L=22nm
Mp9     n7 n2 n5 n5  pmos W=44nm L=22nm
Mp10    n8 a vdd vdd pmos W=44nm L=22nm
Mp11    n9 b n8  n8  pmos W=44nm L=22nm
Mp12    n7 c n9  n9  pmos W=44nm L=22nm

Mp13    n_sum n7 vdd vdd pmos W=44nm L=22nm
Mp14    n_carry n2 vdd vdd pmos W=44nm L=22nm

Mn1     n2 b n1  n1  nmos W=44nm L=22nm
Mn2     n1 a gnd gnd nmos W=44nm L=22nm
Mn3     n2 c n4  n4  nmos W=44nm L=22nm
Mn4     n4 a gnd gnd nmos W=44nm L=22nm
Mn5     n4 b gnd gnd nmos W=44nm L=22nm
Mn6     n6 c gnd gnd nmos W=44nm L=22nm
Mn7     n6 a gnd gnd nmos W=44nm L=22nm
Mn8     n6 b gnd gnd nmos W=44nm L=22nm
Mn9     n7 n2 n6 n6  nmos W=44nm L=22nm
Mn10    n7 c n10 n10 nmos W=44nm L=22nm
Mn11    n10 b n11 n11 nmos W=44nm L=22nm
Mn12    n11 a gnd gnd nmos W=44nm L=22nm

Mn13    n_sum n7 gnd gnd nmos W=44nm L=22nm
Mn14    n_carry n2 gnd gnd nmos W=44nm L=22nm


.ends FullAdder
* ----------------------END OF SUBCIRCUIT----------------------
.end



* -----------------SUBCIRCUIT OF 3-BIT FULL ADDER--------------
.subckt HalfAdder a b n_sum n_carry gnd


Vss3 vdd gnd DC 'SUPPLY'

Mp5 an a vdd vdd pmos W=44nm L=22nm
Mp6 bn b vdd vdd pmos W=44nm L=22nm

Mp1 n_sum b n1 n1 pmos W=44nm L=22nm
Mp2 n_sum bn  n2 n2 pmos W=44nm L=22nm
Mp3 n1 an vdd vdd pmos W=44nm L=22nm
Mp4 n2 a vdd vdd pmos W=44nm L=22nm

Mn5 an a gnd gnd nmos W=44nm L=22nm
Mn6 bn b gnd gnd nmos W=44nm L=22nm

Mn1 n_sum an n3 n3 nmos W=44nm L=22nm
Mn2 n3 bn gnd gnd nmos W=44nm L=22nm
Mn3 n_sum a n4 n4 nmos W=44nm L=22nm
Mn4 n4 b gnd gnd nmos W=44nm L=22nm

* X1 a b n_carry gnd and2


Mp7 nn1 a vdd vdd pmos W=44nm L=22nm
Mp8 nn1 b vdd vdd pmos W=44nm L=22nm
Mp9 n_carry nn1 vdd vdd pmos W=44nm L=22nm

Mn7 nn1 a nn2 nn2 nmos W=44nm L=22nm
Mn8 nn2 b gnd gnd nmos W=44nm L=22nm
Mn9 n_carry nn1 gnd gnd nmos W=44nm L=22nm

.ends HalfAdder
* ----------------------END OF SUBCIRCUIT----------------------
.end




* ----------_INPUT SIGNALS-----------
VinA0 A0 gnd PWL 0ns 0 10ns 0 11ns 'SUPPLY' 20ns 'SUPPLY'
VinA1 A1 gnd PWL 0ns 0 10ns 0 11ns 'SUPPLY' 20ns 'SUPPLY'
VinA2 A2 gnd PWL 0ns 0 10ns 0 11ns 'SUPPLY' 20ns 'SUPPLY'
VinA3 A3 gnd PWL 0ns 0 10ns 0 11ns 'SUPPLY' 20ns 'SUPPLY'

VinB0 B0 gnd PWL 0ns 0 10ns 0 11ns 'SUPPLY' 20ns 'SUPPLY'
VinB1 B1 gnd PWL 0ns 0 10ns 0 11ns 'SUPPLY' 20ns 'SUPPLY'
VinB2 B2 gnd PWL 0ns 0 10ns 0 11ns 'SUPPLY' 20ns 'SUPPLY'
VinB3 B3 gnd PWL 0ns 0 10ns 0 11ns 'SUPPLY' 20ns 'SUPPLY'


* VinA0 A0 gnd 'SUPPLY'
* VinA1 A1 gnd 'SUPPLY'
* VinA2 A2 gnd 'SUPPLY'
* VinA3 A3 gnd 'SUPPLY'

* VinB0 B0 gnd 'SUPPLY'
* VinB1 B1 gnd 'SUPPLY'
* VinB2 B2 gnd 'SUPPLY'
* VinB3 B3 gnd 'SUPPLY'


XHA1  D7  D8  SH1 CH1 gnd HalfAdder
XHA2  S5  C7  P4  CH2 gnd HalfAdder
XHA3  D11 D12 SH3 CH3 gnd HalfAdder
XHA4  D14 D15 P1  PH4 gnd HalfAdder

X1  B3  A3  D1  gnd and2
X2  B2  A3  D2  gnd and2
X3  B3  A2  D3  gnd and2
X4  B3  A1  D4  gnd and2
X5  B1  A3  D5  gnd and2
X6  B2  A2  D6  gnd and2
X7  B1  A2  D7  gnd and2
X8  B0  A3  D8  gnd and2
X9  B3  A0  D9  gnd and2
X10 B2  A1  D10 gnd and2
X11 B1  A1  D11 gnd and2
X12 B0  A2  D12 gnd and2
X13 B2  A0  D13 gnd and2
X14 B0  A1  D14 gnd and2
X15 B1  A0  D15 gnd and2
X16 B0  A0  P0  gnd and2


XFA1 D2  D3  C4  S1  C1  gnd FullAdder
XFA2 D1  C1  C3  P6  C5  gnd FullAdder
XFA3 S1  C5  CH2 P5  C3  gnd FullAdder
XFA4 D5  D6  CH1 S4  C4  gnd FullAdder
XFA5 D4  S4  C6  S5  C5  gnd FullAdder
XFA6 SH1 D10 CH3 S6  C6  gnd FullAdder
XFA7 D9  S6  C8  P3  C7  gnd FullAdder
XFA8 SH3 D13 CH4 P2  C8  gnd FullAdder


.control
tran 10ns 40ns

plot v(A1)
.endc
.end