magic
tech scmos
timestamp 1669307942
<< error_s >>
rect -176 104 -175 107
rect -173 98 -172 104
<< metal1 >>
rect -6491 1037 -6215 1094
rect -6491 950 -6400 1037
rect -6301 950 -6215 1037
rect -6491 872 -6215 950
rect -6025 1015 -5749 1081
rect -6025 928 -5933 1015
rect -5834 928 -5749 1015
rect -6366 523 -6327 872
rect -6025 859 -5749 928
rect -5552 1030 -5276 1087
rect -5552 943 -5464 1030
rect -5365 943 -5276 1030
rect -5552 865 -5276 943
rect -5053 1022 -4777 1087
rect -5053 935 -4969 1022
rect -4870 935 -4777 1022
rect -5053 865 -4777 935
rect -5934 567 -5895 859
rect -5437 606 -5398 865
rect -4940 654 -4901 865
rect -4942 644 -3210 654
rect -4942 643 -799 644
rect -514 643 -481 644
rect -335 643 -302 644
rect -161 643 -128 644
rect -4942 628 -1964 643
rect -1952 629 -18 643
rect -1952 628 -799 629
rect -4942 625 -3210 628
rect -698 627 -665 629
rect -514 628 -481 629
rect -335 628 -302 629
rect -161 628 -128 629
rect -5439 599 -3217 606
rect -700 599 -667 600
rect -5439 589 -2290 599
rect -3241 584 -2290 589
rect -2278 585 -193 599
rect -2278 584 -749 585
rect -700 584 -667 585
rect -3241 583 -749 584
rect -516 583 -483 585
rect -335 583 -302 585
rect -5934 565 -3225 567
rect -5934 558 -2611 565
rect -5926 550 -2611 558
rect -2599 551 -371 565
rect -2599 550 -868 551
rect -5926 549 -868 550
rect -5926 546 -3225 549
rect -6366 522 -3204 523
rect -6366 520 -556 522
rect -6366 507 -2890 520
rect -3241 506 -2890 507
rect -2878 508 -556 520
rect -2878 506 -887 508
rect -1963 330 -1951 332
rect -1964 315 -1963 321
rect -1951 315 -1948 321
rect -1964 306 -1948 315
rect -2278 264 -2277 275
rect -2890 201 -2879 202
rect -2880 186 -2879 201
rect -2890 6 -2879 186
rect -2854 138 -2845 141
rect -2854 128 -2853 138
rect -2846 128 -2845 138
rect -2854 15 -2845 128
rect -2711 22 -2670 26
rect -2854 10 -2837 15
rect -2890 1 -2833 6
rect -2890 -2 -2879 1
rect -2681 -102 -2670 22
rect -2609 8 -2600 211
rect -2568 140 -2560 143
rect -2561 130 -2560 140
rect -2568 17 -2560 130
rect -2534 72 -2527 87
rect -2568 11 -2537 17
rect -2609 2 -2535 8
rect -2409 -88 -2403 28
rect -2289 5 -2277 264
rect -2246 16 -2238 128
rect -2181 72 -2174 87
rect -2078 20 -2030 26
rect -2246 12 -2201 16
rect -2289 -2 -2199 5
rect -2288 -3 -2199 -2
rect -2469 -98 -2403 -88
rect -2782 -115 -2670 -102
rect -2468 -115 -2458 -98
rect -2042 -103 -2031 20
rect -1963 6 -1951 306
rect -1921 15 -1913 128
rect -564 120 -557 508
rect -543 318 -535 324
rect -564 39 -559 120
rect -543 44 -535 303
rect -378 120 -371 551
rect -350 320 -342 323
rect -564 35 -529 39
rect -1751 19 -1691 24
rect -1921 10 -1875 15
rect -1963 1 -1873 6
rect -1963 -1 -1951 1
rect -1724 -94 -1711 19
rect -405 -36 -400 58
rect -378 38 -373 120
rect -350 43 -342 305
rect -200 119 -193 585
rect -183 320 -175 323
rect -183 305 -182 320
rect -378 34 -343 38
rect -977 -41 -397 -36
rect -218 -39 -213 57
rect -199 38 -194 119
rect -183 43 -175 305
rect -25 119 -18 629
rect -4 319 4 322
rect -199 34 -177 38
rect -980 -46 -397 -41
rect -980 -67 -970 -46
rect -219 -64 -213 -39
rect -50 -40 -45 57
rect -24 37 -18 119
rect -4 42 4 304
rect -24 33 3 37
rect 128 -32 133 57
rect -609 -65 -208 -64
rect -2157 -115 -2031 -103
rect -1820 -104 -1711 -94
rect -978 -104 -970 -67
rect -611 -71 -208 -65
rect -611 -78 -603 -71
rect -52 -77 -44 -40
rect -610 -112 -605 -78
rect -294 -85 -40 -77
rect -294 -107 -287 -85
rect -2042 -118 -2031 -115
rect -1820 -739 -1796 -735
rect -3416 -778 -3389 -740
rect -2288 -756 -1795 -739
rect -3416 -801 -2161 -778
rect -4966 -824 -4930 -804
rect -4909 -822 -4883 -804
rect -4909 -824 -2521 -822
rect -4966 -826 -2521 -824
rect -4966 -835 -2516 -826
rect -4966 -838 -4390 -835
rect -4966 -848 -4883 -838
rect -5424 -879 -5419 -852
rect -5390 -861 -5326 -852
rect -5390 -864 -4472 -861
rect -5390 -876 -2936 -864
rect -5390 -879 -4472 -876
rect -5424 -888 -5326 -879
rect -5907 -940 -5879 -914
rect -5850 -917 -5809 -914
rect -5850 -931 -3275 -917
rect -5850 -933 -4511 -931
rect -5850 -940 -5809 -933
rect -5907 -950 -5809 -940
rect -6416 -1002 -6365 -973
rect -6336 -984 -6310 -973
rect -6336 -987 -4754 -984
rect -3700 -987 -3694 -984
rect -6336 -1001 -3691 -987
rect -6336 -1002 -4754 -1001
rect -6416 -1006 -4754 -1002
rect -6416 -1017 -6310 -1006
rect -3700 -1187 -3694 -1001
rect -3654 -1178 -3647 -1065
rect -3510 -1173 -3472 -1168
rect -3654 -1181 -3637 -1178
rect -3700 -1194 -3638 -1187
rect -3493 -1340 -3485 -1173
rect -3291 -1181 -3281 -931
rect -3257 -1173 -3249 -1065
rect -3257 -1176 -3229 -1173
rect -3291 -1188 -3230 -1181
rect -3306 -1332 -3111 -1331
rect -3102 -1332 -3095 -1162
rect -2952 -1178 -2942 -876
rect -2913 -1065 -2912 -1054
rect -2913 -1170 -2904 -1065
rect -2737 -1160 -2733 -1159
rect -2913 -1173 -2866 -1170
rect -2952 -1185 -2866 -1178
rect -2738 -1323 -2733 -1160
rect -2533 -1170 -2516 -835
rect -2504 -1065 -2503 -1054
rect -2494 -1065 -2492 -1054
rect -2504 -1161 -2492 -1065
rect -2504 -1164 -2469 -1161
rect -2504 -1165 -2476 -1164
rect -2533 -1174 -2471 -1170
rect -2346 -1295 -2341 -1152
rect -3602 -1349 -3483 -1340
rect -3306 -1348 -3095 -1332
rect -2968 -1347 -2733 -1323
rect -2617 -1301 -2341 -1295
rect -2617 -1342 -2342 -1301
rect -2737 -1348 -2733 -1347
rect -3290 -1349 -3095 -1348
rect -2192 -1350 -2175 -801
rect -1820 -1346 -1796 -756
rect -1473 -1361 -1439 -742
rect -1128 -767 -813 -731
rect -1126 -1347 -1089 -767
rect -4235 -2038 -4211 -1965
rect -4235 -2040 -3415 -2038
rect -4235 -2059 -3404 -2040
rect -3123 -2042 -3080 -1970
rect -2685 -2021 -2665 -2020
rect -2305 -2021 -2269 -1970
rect -3123 -2047 -3033 -2042
rect -3123 -2056 -3030 -2047
rect -2688 -2050 -2267 -2021
rect -4943 -2161 -3777 -2160
rect -4943 -2183 -4942 -2161
rect -4895 -2183 -3777 -2161
rect -5445 -2253 -5437 -2230
rect -5390 -2253 -4295 -2230
rect -5844 -2305 -4739 -2283
rect -5891 -2306 -4739 -2305
rect -6386 -2380 -6383 -2358
rect -5175 -2358 -5167 -2354
rect -6336 -2380 -5166 -2358
rect -6386 -2381 -5166 -2380
rect -5175 -2588 -5167 -2381
rect -5139 -2579 -5132 -2472
rect -4860 -2568 -4845 -2567
rect -4992 -2575 -4845 -2568
rect -5139 -2584 -5122 -2579
rect -5175 -2595 -5120 -2588
rect -4860 -2791 -4845 -2575
rect -4753 -2576 -4745 -2306
rect -4705 -2566 -4697 -2472
rect -4533 -2563 -4515 -2556
rect -4705 -2572 -4660 -2566
rect -4753 -2581 -4660 -2576
rect -4526 -2796 -4516 -2563
rect -4306 -2568 -4299 -2253
rect -4246 -2474 -4245 -2465
rect -4255 -2557 -4245 -2474
rect -4031 -2547 -4021 -2546
rect -4058 -2554 -4019 -2547
rect -4255 -2561 -4181 -2557
rect -4255 -2563 -4187 -2561
rect -4306 -2573 -4187 -2568
rect -4031 -2783 -4021 -2554
rect -3790 -2568 -3780 -2183
rect -3758 -2558 -3748 -2473
rect -3578 -2554 -3554 -2548
rect -3758 -2562 -3703 -2558
rect -3790 -2574 -3704 -2568
rect -3564 -2778 -3554 -2554
rect -4201 -2800 -4021 -2783
rect -3849 -2792 -3554 -2778
rect -3428 -2793 -3404 -2059
rect -3054 -2800 -3030 -2056
rect -2685 -2788 -2665 -2050
rect -2366 -2090 -2340 -2088
rect -1674 -2090 -1641 -1969
rect -2369 -2126 -1641 -2090
rect -2366 -2788 -2340 -2126
rect -5490 -3890 -5449 -3405
rect -4359 -3890 -4318 -3423
rect -3547 -3890 -3506 -3402
rect -2916 -3890 -2875 -3405
rect -2466 -3890 -2425 -3395
rect -1219 -3890 -1180 -1959
rect -397 -3889 -357 -725
rect 107 -3890 151 -32
rect 396 -90 444 -49
rect 396 -97 399 -90
rect 411 -97 444 -90
rect 396 -669 444 -97
rect 427 -713 444 -669
rect 396 -1243 444 -713
rect 416 -1264 444 -1243
rect 396 -1919 444 -1264
rect 396 -1924 443 -1919
rect 440 -1982 443 -1924
rect 396 -1998 443 -1982
rect 396 -2640 444 -1998
rect 396 -2666 399 -2640
rect 430 -2666 444 -2640
rect 396 -3363 444 -2666
rect 396 -3876 444 -3435
<< m2contact >>
rect -6400 950 -6301 1037
rect -5933 928 -5834 1015
rect -5464 943 -5365 1030
rect -4969 935 -4870 1022
rect -1964 628 -1952 643
rect -2290 584 -2278 599
rect -2611 550 -2599 565
rect -2890 505 -2878 520
rect -1963 315 -1951 330
rect -2290 264 -2278 279
rect -2610 211 -2598 226
rect -2892 186 -2880 201
rect -2853 128 -2846 138
rect -2568 130 -2561 140
rect -2246 128 -2237 135
rect -1921 128 -1913 135
rect -544 303 -535 318
rect -350 305 -341 320
rect -182 305 -173 320
rect -5 304 4 319
rect -4930 -824 -4909 -803
rect -5419 -879 -5390 -849
rect -5879 -940 -5850 -910
rect -6365 -1002 -6336 -972
rect -3656 -1065 -3647 -1051
rect -3257 -1065 -3248 -1054
rect -2912 -1065 -2903 -1054
rect -2503 -1065 -2494 -1054
rect -4942 -2186 -4895 -2161
rect -5437 -2255 -5390 -2230
rect -5891 -2305 -5844 -2280
rect -6383 -2380 -6336 -2355
rect -5140 -2472 -5131 -2463
rect -4705 -2472 -4696 -2463
rect -4255 -2474 -4246 -2465
rect -3758 -2473 -3748 -2460
rect 399 -97 411 -90
rect 394 -713 427 -669
rect 395 -1264 416 -1243
rect 385 -1982 440 -1924
rect 399 -2666 430 -2640
rect 395 -3435 465 -3363
<< metal2 >>
rect -6362 -968 -6337 950
rect -5880 -907 -5860 928
rect -5420 -849 -5398 943
rect -4929 -792 -4909 935
rect -1964 643 -1952 644
rect -2278 584 -2277 598
rect -2610 565 -2597 566
rect -2599 550 -2597 565
rect -2891 520 -2877 524
rect -2891 505 -2890 520
rect -2878 505 -2877 520
rect -3947 158 -3746 219
rect -2891 201 -2877 505
rect -2610 226 -2597 550
rect -2289 279 -2277 584
rect -1964 330 -1952 628
rect -1521 335 -1320 406
rect -1964 315 -1963 330
rect -1521 320 28 335
rect -1521 318 -350 320
rect -1964 314 -1952 315
rect -2278 264 -2277 279
rect -2289 263 -2277 264
rect -1521 303 -544 318
rect -535 305 -350 318
rect -341 305 -182 320
rect -173 319 28 320
rect -173 305 -5 319
rect -535 304 -5 305
rect 4 304 28 319
rect -535 303 28 304
rect -1521 301 28 303
rect -2598 212 -2597 226
rect -1521 210 -1320 301
rect -2880 186 -2877 201
rect -2891 185 -2877 186
rect -3947 140 -1825 158
rect -3947 138 -2568 140
rect -3947 128 -2853 138
rect -2846 130 -2568 138
rect -2561 135 -1825 140
rect -2561 130 -2246 135
rect -2846 128 -2246 130
rect -2237 128 -1921 135
rect -1913 128 -1825 135
rect -3947 127 -1825 128
rect -3947 23 -3746 127
rect 673 122 878 408
rect -2785 116 878 122
rect -2762 76 -2752 116
rect -2477 78 -2467 116
rect -2136 77 -2126 116
rect -1800 75 -1790 116
rect -443 110 -437 116
rect -264 109 -258 116
rect -98 110 -92 116
rect 59 110 65 116
rect -2760 -90 -2751 -28
rect -2504 -90 -2495 -28
rect -2178 -90 -2169 -30
rect -1853 -90 -1844 -28
rect -498 -90 -487 5
rect -255 -90 -244 4
rect -124 -90 -113 4
rect 33 -90 44 3
rect -2795 -97 399 -90
rect 673 -173 878 116
rect 566 -189 878 -173
rect -76 -231 878 -189
rect 566 -232 878 -231
rect -91 -711 394 -669
rect 427 -711 436 -669
rect -4944 -803 -4902 -792
rect -4944 -824 -4930 -803
rect -4909 -824 -4902 -803
rect -5420 -850 -5419 -849
rect -5440 -879 -5419 -850
rect -5390 -879 -5383 -850
rect -5891 -910 -5849 -907
rect -5891 -940 -5879 -910
rect -5850 -940 -5849 -910
rect -6381 -972 -6335 -968
rect -6381 -1002 -6365 -972
rect -6336 -1002 -6335 -972
rect -6381 -2355 -6335 -1002
rect -5891 -2280 -5849 -940
rect -5440 -2230 -5383 -879
rect -4944 -2161 -4902 -824
rect -4506 -1037 -4305 -1026
rect -4506 -1051 -2467 -1037
rect -4506 -1065 -3656 -1051
rect -3647 -1054 -2467 -1051
rect -3647 -1065 -3257 -1054
rect -3248 -1065 -2912 -1054
rect -2903 -1065 -2503 -1054
rect -2494 -1065 -2467 -1054
rect -4506 -1222 -4305 -1065
rect -3585 -1080 -3213 -1078
rect 673 -1080 878 -232
rect -3585 -1092 878 -1080
rect -3585 -1094 -3213 -1092
rect -3567 -1118 -3559 -1094
rect -3187 -1111 -3180 -1092
rect -2813 -1108 -2806 -1092
rect -2401 -1100 -2395 -1092
rect -3563 -1244 -3547 -1221
rect -3164 -1244 -3148 -1216
rect -2829 -1244 -2813 -1215
rect -2426 -1244 -2409 -1203
rect -3563 -1264 395 -1244
rect 416 -1264 444 -1244
rect 673 -1400 878 -1092
rect 553 -1410 878 -1400
rect -948 -1472 878 -1410
rect 553 -1479 878 -1472
rect -1034 -1924 443 -1919
rect -1034 -1981 385 -1924
rect 440 -1981 443 -1924
rect -4944 -2183 -4942 -2161
rect -5440 -2255 -5437 -2230
rect -5390 -2255 -5383 -2230
rect -5891 -2306 -5849 -2305
rect -6336 -2380 -6335 -2355
rect -6381 -2389 -6335 -2380
rect -5501 -2450 -5343 -2411
rect -5501 -2460 -3667 -2450
rect -5501 -2463 -3758 -2460
rect -5501 -2472 -5140 -2463
rect -5131 -2472 -4705 -2463
rect -4696 -2465 -3758 -2463
rect -4696 -2472 -4255 -2465
rect -5501 -2473 -4255 -2472
rect -5501 -2532 -5343 -2473
rect -4246 -2473 -3758 -2465
rect -3748 -2473 -3667 -2460
rect 673 -2482 878 -1479
rect -5222 -2495 878 -2482
rect -5093 -2518 -5082 -2495
rect -4632 -2504 -4624 -2495
rect -5055 -2644 -5050 -2625
rect -4590 -2644 -4585 -2612
rect -4103 -2644 -4097 -2602
rect -3655 -2644 -3649 -2602
rect -5119 -2666 399 -2644
rect 430 -2666 446 -2644
rect 673 -2824 878 -2495
rect -2130 -2924 878 -2824
rect 673 -3047 878 -2924
rect -2166 -3363 533 -3361
rect -2166 -3429 395 -3363
rect 465 -3429 533 -3363
use and  and_7
timestamp 1669290443
transform 1 0 -2837 0 1 -39
box -3 8 130 118
use and  and_6
timestamp 1669290443
transform 1 0 -2537 0 1 -37
box -3 8 130 118
use and  and_5
timestamp 1669290443
transform 1 0 -2200 0 1 -39
box -3 8 130 118
use and  and_4
timestamp 1669290443
transform 1 0 -1875 0 1 -39
box -3 8 130 118
use and  and_3
timestamp 1669290443
transform 1 0 -532 0 1 -6
box -3 8 130 118
use and  and_2
timestamp 1669290443
transform 1 0 -343 0 1 -7
box -3 8 130 118
use and  and_1
timestamp 1669290443
transform 1 0 -177 0 1 -7
box -3 8 130 118
use and  and_0
timestamp 1669290443
transform 1 0 3 0 1 -8
box -3 8 130 118
use 4bitadder  4bitadder_0
timestamp 1669296483
transform 1 0 -432 0 1 -648
box -3434 -106 428 556
use and  and_11
timestamp 1669290443
transform 1 0 -3637 0 1 -1232
box -3 8 130 118
use and  and_10
timestamp 1669290443
transform 1 0 -3229 0 1 -1227
box -3 8 130 118
use and  and_9
timestamp 1669290443
transform 1 0 -2866 0 1 -1224
box -3 8 130 118
use and  and_8
timestamp 1669290443
transform 1 0 -2473 0 1 -1215
box -3 8 130 118
use 4bitadder  4bitadder_1
timestamp 1669296483
transform 1 0 -1255 0 1 -1885
box -3434 -106 428 556
use and  and_12
timestamp 1669290443
transform 1 0 -5119 0 1 -2634
box -3 8 130 118
use and  and_13
timestamp 1669290443
transform 1 0 -4659 0 1 -2621
box -3 8 130 118
use and  and_14
timestamp 1669290443
transform 1 0 -4186 0 1 -2612
box -3 8 130 118
use and  and_15
timestamp 1669290443
transform 1 0 -3704 0 1 -2612
box -3 8 130 118
use 4bitadder  4bitadder_2
timestamp 1669296483
transform 1 0 -2495 0 1 -3330
box -3434 -106 428 556
<< end >>
