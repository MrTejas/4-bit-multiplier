* SPICE3 file created from inverter_test.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY=5
.option scale=0.09u
.global vdd gnd


Vdd vdd gnd 'SUPPLY'
vinA input gnd pulse 0 'SUPPLY' 0ns 0.5ns 0.5ns 10ns 20ns


M1000 out1 input gnd Gnd nfet w=4 l=2
+  ad=20 pd=18 as=20 ps=18
M1001 out1 input vdd inverter_0/w_0_0# pfet w=9 l=2
+  ad=45 pd=28 as=54 ps=30
C0 vdd out1 0.10fF
C1 inverter_0/w_0_0# vdd 0.10fF
C2 inverter_0/w_0_0# out1 0.04fF
C3 input out1 0.03fF
C4 out1 gnd 0.07fF
C5 inverter_0/w_0_0# input 0.08fF
C6 input gnd 0.02fF
C7 gnd Gnd 0.14fF
C8 out1 Gnd 0.15fF
C9 vdd Gnd 0.05fF
C10 input Gnd 0.24fF
C11 inverter_0/w_0_0# Gnd 0.73fF




.tran 0.1n 40n

.control
* set hcopycolor = 1
* set color0=white
* set color1=black

run
plot v(input) v(out1)+6

.endc

.end