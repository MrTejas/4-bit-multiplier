magic
tech scmos
timestamp 1669308879
<< error_s >>
rect 6317 3995 6318 3998
rect 6320 3989 6321 3995
<< metal1 >>
rect 84 4937 208 5022
rect 597 4925 721 5010
rect 1028 4936 1152 5021
rect 1523 4926 1647 5011
rect 5118 3801 5144 3812
rect 5118 3794 5122 3801
rect 5135 3794 5144 3801
rect 5118 3792 5144 3794
rect 958 -27 1082 58
rect 2075 -14 2199 71
rect 2891 -22 3015 63
rect 3547 -2 3671 83
rect 3987 -5 4111 80
rect 5216 -7 5340 78
rect 6038 5 6162 90
rect 6551 -1 6675 84
rect 6869 16 6993 101
<< m2contact >>
rect 5122 3794 5135 3801
<< metal2 >>
rect 5024 4138 5148 4223
rect 7101 4151 7424 4363
rect 2589 3954 2713 4039
rect 2026 2714 2150 2799
rect 1009 1385 1133 1470
use multiplier  multiplier_0
timestamp 1669307942
transform 1 0 6493 0 1 3891
box -6491 -3890 878 1094
<< labels >>
rlabel metal1 102 4942 168 4984 1 inA3
rlabel metal1 618 4931 684 4973 1 inA2
rlabel metal1 1048 4937 1114 4979 1 inA1
rlabel metal1 1551 4936 1617 4978 1 inA0
rlabel metal2 5043 4160 5109 4202 1 inB0
rlabel metal2 2617 3972 2683 4014 1 inB1
rlabel metal2 2057 2728 2123 2770 1 inB2
rlabel metal2 1028 1395 1094 1437 1 inB3
rlabel metal1 6601 9 6639 54 1 P0
rlabel metal1 6100 17 6138 62 1 P1
rlabel metal1 5268 14 5306 59 1 P2
rlabel metal1 4033 22 4071 67 1 P3
rlabel metal1 3581 14 3619 59 1 P4
rlabel metal1 2948 10 2986 55 1 P5
rlabel metal1 2131 7 2169 52 1 P6
rlabel metal1 1004 1 1042 46 1 P7
rlabel metal1 6891 30 6924 63 1 gnd
rlabel metal2 7215 4214 7262 4277 1 vdd
<< end >>
