magic
tech scmos
timestamp 1669296483
<< metal1 >>
rect -2373 521 -2331 541
rect -2373 508 -2362 521
rect -2348 508 -2331 521
rect -2065 520 -2023 539
rect -2065 507 -2049 520
rect -2036 507 -2023 520
rect -1730 522 -1688 543
rect -1730 510 -1716 522
rect -1704 510 -1688 522
rect -1387 527 -1345 549
rect -1387 516 -1372 527
rect -1362 516 -1345 527
rect -948 519 -904 552
rect -567 522 -523 555
rect -198 523 -154 556
rect 119 523 163 556
rect -2065 506 -2023 507
rect -934 494 -913 519
rect -2964 485 -913 494
rect -3091 379 -3083 466
rect -2964 384 -2956 485
rect -557 479 -539 522
rect -1833 472 -539 479
rect -2858 385 -2249 398
rect -3416 206 -3377 215
rect -3416 17 -3404 206
rect -2264 202 -2250 385
rect -1960 376 -1952 463
rect -1832 379 -1824 472
rect -557 471 -539 472
rect -186 468 -172 523
rect -1726 385 -1125 398
rect -1134 213 -1126 385
rect -827 381 -816 461
rect -698 463 -172 468
rect -698 381 -687 463
rect -594 383 3 391
rect -1134 205 -1119 213
rect -4 112 3 383
rect 129 261 134 473
rect 139 261 143 523
rect 412 128 427 139
rect -3416 -5 -2953 17
rect -2255 12 -1823 13
rect -2981 -92 -2953 -5
rect -2898 -6 -1823 12
rect -634 6 -390 7
rect -2255 -7 -1823 -6
rect -1859 -104 -1825 -7
rect -1766 -11 -1014 5
rect -634 -10 -386 6
rect -1046 -106 -1014 -11
rect -413 -98 -386 -10
rect 36 -8 54 -7
rect 415 -8 427 128
rect 36 -16 428 -8
rect 36 -89 54 -16
<< m2contact >>
rect -2362 508 -2348 521
rect -2049 507 -2036 520
rect -1716 510 -1704 522
rect -1372 516 -1362 527
rect -3092 466 -3083 478
rect -1960 463 -1952 474
rect 125 473 134 483
rect -827 461 -816 468
<< metal2 >>
rect -2362 478 -2348 508
rect -3083 466 -2348 478
rect -2049 474 -2036 507
rect -2049 463 -1960 474
rect -1716 468 -1704 510
rect -1372 483 -1362 516
rect -1372 473 125 483
rect -1716 461 -827 468
rect -931 454 -917 455
rect -3434 422 413 454
rect -3179 359 -3164 422
rect -2040 360 -2025 422
rect -931 359 -917 422
rect 199 251 214 422
rect -3122 -22 -3107 54
rect -2053 -22 -2038 51
rect -895 -22 -881 57
rect 285 -22 297 5
rect -3434 -54 413 -22
use fulladder  fulladder_2
timestamp 1669293643
transform 1 0 -3218 0 1 82
box -168 -81 938 308
use fulladder  fulladder_1
timestamp 1669293643
transform 1 0 -2087 0 1 79
box -168 -81 938 308
use fulladder  fulladder_0
timestamp 1669293643
transform 1 0 -954 0 1 81
box -168 -81 938 308
use halfadder  halfadder_0
timestamp 1669290883
transform 1 0 174 0 1 5
box -174 -5 241 260
<< end >>
